//: version "1.8.7"

module CaLoA(cf, p, g, ci);
//: interface  /sz:(40, 40) /bd:[ Ti0>p(10/40) Ti1>g(28/40) Ri0>ci(22/40) Lo0<cf(20/40) ]
input p;    //: /sn:0 {0}(105,123)(163,123)(163,134)(173,134){1}
output cf;    //: /sn:0 /dp:1 {0}(261,99)(319,99){1}
input ci;    //: /sn:0 {0}(109,150)(163,150)(163,139)(173,139){1}
input g;    //: /sn:0 {0}(107,87)(230,87)(230,96)(240,96){1}
wire w2;    //: /sn:0 {0}(194,137)(230,137)(230,101)(240,101){1}
//: enddecls

  xor g4 (.I0(p), .I1(ci), .Z(w2));   //: @(184,137) /sn:0 /w:[ 1 1 0 ]
  //: output g3 (cf) @(316,99) /sn:0 /w:[ 1 ]
  //: input g2 (p) @(103,123) /sn:0 /w:[ 0 ]
  //: input g1 (g) @(105,87) /sn:0 /w:[ 0 ]
  and g5 (.I0(g), .I1(w2), .Z(cf));   //: @(251,99) /sn:0 /w:[ 1 1 0 ]
  //: input g0 (ci) @(107,150) /sn:0 /w:[ 0 ]

endmodule

module Carrylookahead_logic(p3, g3, c3, c2, c1, p1, g0, c4, g2, g1, p2, c0, p0);
//: interface  /sz:(379, 40) /bd:[ Ti0>g0(321/379) Ti1>p0(311/379) Ti2>g1(233/379) Ti3>p1(225/379) Ti4>g2(144/379) Ti5>p2(135/379) Ti6>g3(58/379) Ti7>p3(50/379) Ri0>c0(24/40) To0<c3(95/379) To1<c2(182/379) To2<c1(272/379) Lo0<c4(20/40) ]
input g3;    //: /sn:0 {0}(179,35)(179,120){1}
input g2;    //: /sn:0 {0}(243,35)(243,82)(242,82)(242,122){1}
input g1;    //: /sn:0 {0}(327,35)(327,88)(329,88)(329,124){1}
input c0;    //: /sn:0 {0}(64,-33)(509,-33)(509,149)(441,149){1}
output c1;    //: /sn:0 {0}(38,-16)(379,-16)(379,145){1}
//: {2}(381,147)(399,147){3}
//: {4}(377,147)(360,147){5}
output c4;    //: /sn:0 {0}(150,141)(30,141){1}
input p3;    //: /sn:0 {0}(158,35)(158,82)(161,82)(161,120){1}
input p2;    //: /sn:0 {0}(260,35)(260,122){1}
input p1;    //: /sn:0 {0}(343,34)(343,87)(347,87)(347,124){1}
output c3;    //: /sn:0 {0}(38,15)(209,15)(209,141){1}
//: {2}(211,143)(231,143){3}
//: {4}(207,143)(192,143){5}
input p0;    //: /sn:0 {0}(412,41)(412,90)(410,90)(410,126){1}
output c2;    //: /sn:0 {0}(69,0)(298,0)(298,143){1}
//: {2}(300,145)(318,145){3}
//: {4}(296,145)(273,145){5}
input g0;    //: /sn:0 {0}(429,40)(429,94)(428,94)(428,126){1}
//: enddecls

  //: input g8 (p3) @(158,33) /sn:0 /R:3 /w:[ 0 ]
  CaLoA g4 (.g(g3), .p(p3), .ci(c3), .cf(c4));   //: @(151, 121) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<0 ]
  //: input g13 (g3) @(179,33) /sn:0 /R:3 /w:[ 0 ]
  //: output g3 (c3) @(41,15) /sn:0 /R:2 /w:[ 0 ]
  //: output g2 (c2) @(72,0) /sn:0 /R:2 /w:[ 0 ]
  //: output g1 (c1) @(41,-16) /sn:0 /R:2 /w:[ 0 ]
  //: input g16 (p1) @(343,32) /sn:0 /R:3 /w:[ 0 ]
  //: joint g11 (c2) @(298, 145) /w:[ 2 1 4 -1 ]
  //: joint g10 (c1) @(379, 147) /w:[ 2 1 4 -1 ]
  //: input g19 (g0) @(429,38) /sn:0 /R:3 /w:[ 0 ]
  CaLoA g6 (.g(p1), .p(g1), .ci(c1), .cf(c2));   //: @(319, 125) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<3 ]
  //: output g9 (c4) @(33,141) /sn:0 /R:2 /w:[ 1 ]
  CaLoA g7 (.g(g0), .p(p0), .ci(c0), .cf(c1));   //: @(400, 127) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<3 ]
  //: input g15 (g2) @(243,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g17 (g1) @(327,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g14 (p2) @(260,33) /sn:0 /R:3 /w:[ 0 ]
  CaLoA g5 (.g(p2), .p(g2), .ci(c2), .cf(c3));   //: @(232, 123) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<3 ]
  //: input g0 (c0) @(62,-33) /sn:0 /w:[ 0 ]
  //: input g18 (p0) @(412,39) /sn:0 /R:3 /w:[ 0 ]
  //: joint g12 (c3) @(209, 143) /w:[ 2 1 4 -1 ]

endmodule

module main;    //: root_module
supply0 w20;    //: /sn:0 {0}(685,212)(685,202)(645,202)(645,261)(651,261){1}
wire w32;    //: /sn:0 {0}(522,427)(522,333){1}
//: {2}(524,331)(651,331){3}
//: {4}(520,331)(492,331)(492,110){5}
wire w6;    //: /sn:0 /dp:1 {0}(101,65)(101,18){1}
//: {2}(103,16)(150,16)(150,11){3}
//: {4}(101,14)(101,-23){5}
wire w7;    //: /sn:0 /dp:1 {0}(-76,64)(-76,42){1}
//: {2}(-74,40)(-27,40)(-27,32){3}
//: {4}(-76,38)(-76,-23){5}
wire w61;    //: /sn:0 {0}(560,-71)(560,13){1}
//: {2}(562,15)(591,15)(591,2){3}
//: {4}(560,17)(560,76){5}
wire w46;    //: /sn:0 /dp:1 {0}(290,115)(290,196)(294,196)(294,198){1}
wire w14;    //: /sn:0 {0}(486,-23)(486,39){1}
//: {2}(488,41)(529,41)(529,30){3}
//: {4}(486,43)(486,68){5}
wire w16;    //: /sn:0 {0}(675,96)(638,96){1}
//: {2}(634,96)(587,96){3}
//: {4}(636,98)(636,223)(624,223){5}
wire w4;    //: /sn:0 /dp:1 {0}(0,64)(0,14){1}
//: {2}(2,12)(38,12)(38,-6){3}
//: {4}(0,10)(0,-71){5}
wire w38;    //: /sn:0 {0}(-2,106)(-2,184)(2,184)(2,194){1}
wire w3;    //: /sn:0 {0}(-41,194)(-41,129)(-47,129)(-47,84)(-62,84){1}
wire w0;    //: /sn:0 /dp:1 {0}(-175,64)(-175,34){1}
//: {2}(-173,32)(-123,32)(-123,26){3}
//: {4}(-175,30)(-175,-71){5}
wire w64;    //: /sn:0 {0}(558,118)(558,188)(555,188)(555,198){1}
wire w37;    //: /sn:0 {0}(426,198)(426,89)(408,89){1}
wire w34;    //: /sn:0 {0}(339,198)(339,93)(319,93){1}
wire w21;    //: /sn:0 {0}(-144,415)(-144,390)(-133,390)(-133,273){1}
//: {2}(-131,271)(651,271){3}
//: {4}(-135,271)(-158,271)(-158,106){5}
wire w43;    //: /sn:0 {0}(243,219)(228,219)(228,163){1}
//: {2}(228,159)(228,122){3}
//: {4}(226,161)(197,161)(197,165)(191,165){5}
//: {6}(189,163)(189,85)(115,85){7}
//: {8}(189,167)(189,219)(157,219){9}
wire w31;    //: /sn:0 {0}(440,420)(440,379)(437,379)(437,323){1}
//: {2}(439,321)(651,321){3}
//: {4}(435,321)(398,321)(398,111){5}
wire w58;    //: /sn:0 {0}(471,110)(471,183)(469,183)(469,198){1}
wire w28;    //: /sn:0 {0}(171,419)(171,373)(170,373)(170,293){1}
//: {2}(172,291)(651,291){3}
//: {4}(168,291)(17,291)(17,106){5}
wire [7:0] w24;    //: /sn:0 /dp:8 {0}(-273,-75)(-176,-75){1}
//: {2}(-175,-75)(-90,-75){3}
//: {4}(-89,-75)(-1,-75){5}
//: {6}(0,-75)(87,-75){7}
//: {8}(88,-75)(291,-75){9}
//: {10}(292,-75)(380,-75){11}
//: {12}(381,-75)(474,-75){13}
//: {14}(475,-75)(559,-75){15}
//: {16}(560,-75)(638,-75){17}
wire w41;    //: /sn:0 {0}(86,107)(86,184)(88,184)(88,194){1}
wire w36;    //: /sn:0 {0}(-81,106)(-81,184)(-79,184)(-79,194){1}
wire w1;    //: /sn:0 /dp:1 {0}(-162,64)(-162,50){1}
//: {2}(-160,48)(-110,48)(-110,42){3}
//: {4}(-162,46)(-162,-23){5}
wire [7:0] w25;    //: /sn:0 /dp:8 {0}(-275,-27)(-163,-27){1}
//: {2}(-162,-27)(-77,-27){3}
//: {4}(-76,-27)(12,-27){5}
//: {6}(13,-27)(100,-27){7}
//: {8}(101,-27)(304,-27){9}
//: {10}(305,-27)(393,-27){11}
//: {12}(394,-27)(485,-27){13}
//: {14}(486,-27)(572,-27){15}
//: {16}(573,-27)(634,-27){17}
wire w65;    //: /sn:0 {0}(568,118)(568,188)(565,188)(565,198){1}
wire w40;    //: /sn:0 {0}(516,198)(516,88)(502,88){1}
wire w8;    //: /sn:0 {0}(-165,194)(-165,135)(-167,135)(-167,106){1}
wire w35;    //: /sn:0 {0}(-91,106)(-91,184)(-88,184)(-88,194){1}
wire w18;    //: /sn:0 {0}(88,-71)(88,-4){1}
//: {2}(90,-2)(139,-2)(139,-10){3}
//: {4}(88,0)(88,65){5}
wire w30;    //: /sn:0 {0}(351,425)(351,366)(346,366)(346,313){1}
//: {2}(348,311)(651,311){3}
//: {4}(344,311)(309,311)(309,115){5}
wire w22;    //: /sn:0 {0}(-39,420)(-39,356)(-41,356)(-41,283){1}
//: {2}(-39,281)(57,281){3}
//: {4}(61,281)(651,281){5}
//: {6}(59,283)(59,418){7}
//: {8}(-43,281)(-72,281)(-72,106){9}
wire w17;    //: /sn:0 {0}(-238,126)(-238,215)(-224,215){1}
wire w59;    //: /sn:0 {0}(483,110)(483,190)(477,190)(477,198){1}
wire w53;    //: /sn:0 {0}(389,111)(389,186)(388,186)(388,198){1}
wire w62;    //: /sn:0 {0}(573,-23)(573,31){1}
//: {2}(575,33)(606,33)(606,27){3}
//: {4}(573,35)(573,76){5}
wire w49;    //: /sn:0 {0}(381,-71)(381,28){1}
//: {2}(383,30)(428,30)(428,10){3}
//: {4}(381,32)(381,69){5}
wire w44;    //: /sn:0 {0}(305,-23)(305,25){1}
//: {2}(307,27)(344,27)(344,17){3}
//: {4}(305,29)(305,73){5}
wire w2;    //: /sn:0 {0}(-128,194)(-128,84)(-148,84){1}
wire w11;    //: /sn:0 {0}(-89,64)(-89,19){1}
//: {2}(-87,17)(-47,17)(-47,7){3}
//: {4}(-89,15)(-89,-71){5}
wire [8:0] w10;    //: /sn:0 /dp:1 {0}(768,301)(657,301){1}
wire w13;    //: /sn:0 {0}(13,-23)(13,29){1}
//: {2}(15,31)(51,31)(51,18){3}
//: {4}(13,33)(13,64){5}
wire w33;    //: /sn:0 {0}(606,421)(606,383)(602,383)(602,343){1}
//: {2}(604,341)(651,341){3}
//: {4}(600,341)(577,341)(577,118){5}
wire w52;    //: /sn:0 {0}(379,111)(379,198){1}
wire w5;    //: /sn:0 {0}(49,194)(49,132)(43,132)(43,84)(27,84){1}
wire w29;    //: /sn:0 {0}(279,426)(279,357)(272,357)(272,303){1}
//: {2}(274,301)(651,301){3}
//: {4}(270,301)(105,301)(105,107){5}
wire w47;    //: /sn:0 /dp:1 {0}(300,115)(300,188)(302,188)(302,198){1}
wire w50;    //: /sn:0 {0}(394,-23)(394,42){1}
//: {2}(396,44)(439,44)(439,32){3}
//: {4}(394,46)(394,69){5}
wire w9;    //: /sn:0 {0}(-173,194)(-173,134)(-177,134)(-177,106){1}
wire w42;    //: /sn:0 {0}(96,107)(96,184)(98,184)(98,194){1}
wire w55;    //: /sn:0 {0}(475,-71)(475,24){1}
//: {2}(477,26)(515,26)(515,6){3}
//: {4}(475,28)(475,68){5}
wire w26;    //: /sn:0 {0}(292,-71)(292,8){1}
//: {2}(294,10)(329,10)(329,-2){3}
//: {4}(292,12)(292,73){5}
wire w39;    //: /sn:0 {0}(8,106)(8,184)(10,184)(10,194){1}
//: enddecls

  //: dip g4 (w24) @(-311,-75) /sn:0 /R:1 /w:[ 0 ] /st:22
  tran g8(.Z(w4), .I(w24[5]));   //: @(0,-77) /sn:0 /R:1 /w:[ 5 5 6 ] /ss:1
  led g61 (.I(w1));   //: @(-110,35) /sn:0 /w:[ 3 ] /type:0
  led g51 (.I(w32));   //: @(522,434) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g37 (w22) @(59, 281) /w:[ 4 -1 3 6 ]
  //: supply0 g34 (w20) @(685,218) /sn:0 /w:[ 0 ]
  S_CLA g3 (.B(w6), .A(w18), .C(w43), .S(w29), .G(w42), .P(w41));   //: @(74, 66) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>5 Ri0>7 Bo0<5 Bo1<0 Bo2<0 ]
  tran g13(.Z(w1), .I(w25[7]));   //: @(-162,-29) /sn:0 /R:1 /w:[ 5 1 2 ] /ss:1
  led g58 (.I(w18));   //: @(139,-17) /sn:0 /w:[ 3 ] /type:0
  //: joint g55 (w0) @(-175, 32) /w:[ 2 4 -1 1 ]
  S_CLA g2 (.B(w13), .A(w4), .C(w5), .S(w28), .G(w39), .P(w38));   //: @(-14, 65) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>0 Ri0>1 Bo0<5 Bo1<0 Bo2<0 ]
  //: joint g65 (w18) @(88, -2) /w:[ 2 1 -1 4 ]
  led g76 (.I(w14));   //: @(529,23) /sn:0 /w:[ 3 ] /type:0
  led g77 (.I(w62));   //: @(606,20) /sn:0 /w:[ 3 ] /type:0
  led g59 (.I(w7));   //: @(-27,25) /sn:0 /w:[ 3 ] /type:0
  S_CLA g1 (.B(w7), .A(w11), .C(w3), .S(w22), .G(w36), .P(w35));   //: @(-103, 65) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<9 Bo1<0 Bo2<0 ]
  //: joint g72 (w26) @(292, 10) /w:[ 2 1 -1 4 ]
  led g64 (.I(w26));   //: @(329,-9) /sn:0 /w:[ 3 ] /type:0
  tran g11(.Z(w6), .I(w25[4]));   //: @(101,-29) /sn:0 /R:1 /w:[ 5 7 8 ] /ss:1
  Carrylookahead_logic g16 (.p3(w9), .g3(w8), .p2(w35), .g2(w36), .p1(w38), .g1(w39), .p0(w41), .g0(w42), .c0(w43), .c1(w5), .c2(w3), .c3(w2), .c4(w17));   //: @(-223, 195) /sz:(379, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>9 To0<0 To1<0 To2<0 Lo0<1 ]
  //: joint g87 (w43) @(228, 161) /w:[ -1 2 4 1 ]
  led g50 (.I(w31));   //: @(440,427) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g28 (.I(w17));   //: @(-238,119) /sn:0 /w:[ 0 ] /type:0
  tran g10(.Z(w13), .I(w25[5]));   //: @(13,-29) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  led g78 (.I(w61));   //: @(591,-5) /sn:0 /w:[ 3 ] /type:0
  tran g27(.Z(w62), .I(w25[0]));   //: @(573,-29) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  S_CLA g19 (.B(w50), .A(w49), .C(w37), .S(w31), .G(w53), .P(w52));   //: @(367, 70) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<5 Bo1<0 Bo2<0 ]
  led g32 (.I(w10));   //: @(775,301) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: joint g38 (w28) @(170, 291) /w:[ 2 -1 4 1 ]
  tran g6(.Z(w0), .I(w24[7]));   //: @(-175,-77) /sn:0 /R:1 /w:[ 5 1 2 ] /ss:1
  //: joint g69 (w1) @(-162, 48) /w:[ 2 4 -1 1 ]
  tran g7(.Z(w11), .I(w24[6]));   //: @(-89,-77) /sn:0 /R:1 /w:[ 5 3 4 ] /ss:1
  tran g9(.Z(w18), .I(w24[4]));   //: @(88,-77) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  led g57 (.I(w13));   //: @(51,11) /sn:0 /w:[ 3 ] /type:0
  led g53 (.I(w49));   //: @(428,3) /sn:0 /w:[ 3 ] /type:0
  led g75 (.I(w55));   //: @(515,-1) /sn:0 /w:[ 3 ] /type:0
  tran g31(.Z(w44), .I(w25[3]));   //: @(305,-29) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  S_CLA g20 (.B(w14), .A(w55), .C(w40), .S(w32), .G(w59), .P(w58));   //: @(461, 69) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<5 Bo1<0 Bo2<0 ]
  Carrylookahead_logic g15 (.p3(w46), .g3(w47), .p2(w52), .g2(w53), .p1(w58), .g1(w59), .p0(w64), .g0(w65), .c0(w16), .c1(w40), .c2(w37), .c3(w34), .c4(w43));   //: @(244, 199) /sz:(379, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<0 ]
  //: joint g71 (w7) @(-76, 40) /w:[ 2 4 -1 1 ]
  //: joint g39 (w29) @(272, 301) /w:[ 2 -1 4 1 ]
  //: joint g67 (w13) @(13, 31) /w:[ 2 1 -1 4 ]
  //: joint g68 (w4) @(0, 12) /w:[ 2 4 -1 1 ]
  led g48 (.I(w29));   //: @(279,433) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g43 (w33) @(602, 341) /w:[ 2 -1 4 1 ]
  //: joint g88 (w43) @(189, 165) /w:[ 5 6 -1 8 ]
  tran g29(.Z(w50), .I(w25[2]));   //: @(394,-29) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  tran g25(.Z(w55), .I(w24[1]));   //: @(475,-77) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  led g62 (.I(w6));   //: @(150,4) /sn:0 /w:[ 3 ] /type:0
  //: joint g73 (w44) @(305, 27) /w:[ 2 1 -1 4 ]
  led g17 (.I(w43));   //: @(228,115) /sn:0 /w:[ 3 ] /type:0
  led g52 (.I(w33));   //: @(606,428) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g42 (w32) @(522, 331) /w:[ 2 -1 4 1 ]
  led g63 (.I(w44));   //: @(344,10) /sn:0 /w:[ 3 ] /type:0
  //: joint g83 (w50) @(394, 44) /w:[ 2 1 -1 4 ]
  led g74 (.I(w50));   //: @(439,25) /sn:0 /w:[ 3 ] /type:0
  //: dip g5 (w25) @(-313,-27) /sn:0 /R:1 /w:[ 0 ] /st:22
  //: switch g14 (w16) @(693,96) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g56 (.I(w4));   //: @(38,-13) /sn:0 /w:[ 3 ] /type:0
  led g47 (.I(w28));   //: @(171,426) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g44 (.I(w21));   //: @(-144,422) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g79 (w62) @(573, 33) /w:[ 2 1 -1 4 ]
  //: joint g80 (w61) @(560, 15) /w:[ 2 1 -1 4 ]
  //: joint g36 (w22) @(-41, 281) /w:[ 2 -1 8 1 ]
  tran g24(.Z(w49), .I(w24[2]));   //: @(381,-77) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  S_CLA g21 (.B(w62), .A(w61), .C(w16), .S(w33), .G(w65), .P(w64));   //: @(546, 77) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>3 Bo0<5 Bo1<0 Bo2<0 ]
  //: joint g84 (w49) @(381, 30) /w:[ 2 1 -1 4 ]
  //: joint g41 (w31) @(437, 321) /w:[ 2 -1 4 1 ]
  tran g23(.Z(w26), .I(w24[3]));   //: @(292,-77) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: joint g40 (w30) @(346, 311) /w:[ 2 -1 4 1 ]
  led g54 (.I(w0));   //: @(-123,19) /sn:0 /w:[ 3 ] /type:0
  led g60 (.I(w11));   //: @(-47,0) /sn:0 /w:[ 3 ] /type:0
  //: joint g81 (w14) @(486, 41) /w:[ 2 1 -1 4 ]
  led g46 (.I(w22));   //: @(59,425) /sn:0 /R:2 /w:[ 7 ] /type:0
  led g45 (.I(w22));   //: @(-39,427) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: joint g35 (w21) @(-133, 271) /w:[ 2 -1 4 1 ]
  tran g26(.Z(w61), .I(w24[0]));   //: @(560,-77) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: joint g22 (w16) @(636, 96) /w:[ 1 -1 2 4 ]
  S_CLA g0 (.B(w1), .A(w0), .C(w2), .S(w21), .G(w8), .P(w9));   //: @(-189, 65) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<5 Bo1<1 Bo2<1 ]
  //: joint g70 (w11) @(-89, 17) /w:[ 2 4 -1 1 ]
  //: joint g66 (w6) @(101, 16) /w:[ 2 4 -1 1 ]
  //: joint g82 (w55) @(475, 26) /w:[ 2 1 -1 4 ]
  S_CLA g18 (.B(w44), .A(w26), .C(w34), .S(w30), .G(w47), .P(w46));   //: @(278, 74) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Bo0<5 Bo1<0 Bo2<0 ]
  tran g12(.Z(w7), .I(w25[6]));   //: @(-76,-29) /sn:0 /R:1 /w:[ 5 3 4 ] /ss:1
  tran g33(.Z(w14), .I(w25[1]));   //: @(486,-29) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  concat g30 (.I0(w33), .I1(w32), .I2(w31), .I3(w30), .I4(w29), .I5(w28), .I6(w22), .I7(w21), .I8(w20), .Z(w10));   //: @(656,301) /sn:0 /w:[ 3 3 3 3 3 3 5 3 1 1 ] /dr:0
  led g49 (.I(w30));   //: @(351,432) /sn:0 /R:2 /w:[ 0 ] /type:0

endmodule

module S_CLA(P, A, C, G, S, B);
//: interface  /sz:(40, 40) /bd:[ Ti0>A(14/40) Ti1>B(27/40) Ri0>C(19/40) Bo0<P(12/40) Bo1<G(22/40) Bo2<S(31/40) ]
input B;    //: /sn:0 {0}(-293,-95)(-250,-95){1}
//: {2}(-246,-95)(-223,-95)(-223,-105)(-149,-105){3}
//: {4}(-248,-93)(-248,-74){5}
//: {6}(-246,-72)(-35,-72){7}
//: {8}(-248,-70)(-248,-34)(-36,-34){9}
input A;    //: /sn:0 /dp:1 {0}(-149,-110)(-222,-110)(-222,-119)(-269,-119){1}
//: {2}(-273,-119)(-294,-119){3}
//: {4}(-271,-117)(-271,-69){5}
//: {6}(-269,-67)(-35,-67){7}
//: {8}(-271,-65)(-271,-29)(-36,-29){9}
output G;    //: /sn:0 /dp:1 {0}(-15,-31)(73,-31){1}
input C;    //: /sn:0 {0}(-293,-80)(-62,-80)(-62,-120)(-37,-120){1}
output P;    //: /sn:0 {0}(73,-69)(-14,-69){1}
output S;    //: /sn:0 /dp:1 {0}(-16,-122)(73,-122){1}
wire w3;    //: /sn:0 /dp:1 {0}(-37,-125)(-76,-125)(-76,-107)(-128,-107){1}
//: enddecls

  //: output g8 (P) @(70,-69) /sn:0 /w:[ 0 ]
  //: input g4 (A) @(-296,-119) /sn:0 /w:[ 3 ]
  //: joint g13 (B) @(-248, -72) /w:[ 6 5 -1 8 ]
  and g3 (.I0(B), .I1(A), .Z(G));   //: @(-25,-31) /sn:0 /w:[ 9 9 0 ]
  or g2 (.I0(B), .I1(A), .Z(P));   //: @(-24,-69) /sn:0 /w:[ 7 7 1 ]
  xor g1 (.I0(w3), .I1(C), .Z(S));   //: @(-26,-122) /sn:0 /w:[ 0 1 0 ]
  //: joint g11 (A) @(-271, -67) /w:[ 6 5 -1 8 ]
  //: joint g10 (A) @(-271, -119) /w:[ 1 -1 2 4 ]
  //: input g6 (C) @(-295,-80) /sn:0 /w:[ 0 ]
  //: output g9 (G) @(70,-31) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(70,-122) /sn:0 /w:[ 1 ]
  //: input g5 (B) @(-295,-95) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(w3));   //: @(-138,-107) /sn:0 /w:[ 0 3 1 ]
  //: joint g12 (B) @(-248, -95) /w:[ 2 -1 1 4 ]

endmodule
