//: version "1.8.7"

module Data_Memory(WriteData, MemWrite, Address, MemRead, ReadData);
//: interface  /sz:(117, 144) /bd:[ Ti0>MemWrite(73/117) Ti1>MemWrite(73/117) Li0>WriteData[31:0](96/144) Li1>Address[31:0](44/144) Li2>WriteData[31:0](96/144) Li3>Address[31:0](44/144) Bi0>MemRead(65/117) Bi1>MemRead(65/117) Ro0<ReadData[31:0](84/144) Ro1<ReadData[31:0](84/144) ]
supply0 w1;    //: /sn:0 {0}(202,264)(202,225){1}
input MemWrite;    //: /sn:0 {0}(151,111)(209,111)(209,122){1}
//: {2}(211,124)(261,124)(261,135){3}
//: {4}(209,126)(209,175){5}
input [31:0] Address;    //: /sn:0 {0}(88,213)(135,213)(135,200){1}
//: {2}(135,199)(135,190){3}
output [31:0] ReadData;    //: /sn:0 {0}(269,140)(277,140)(277,196){1}
//: {2}(279,198)(306,198){3}
//: {4}(275,198)(226,198){5}
input [31:0] WriteData;    //: /sn:0 {0}(193,82)(243,82)(243,140)(253,140){1}
input MemRead;    //: /sn:0 {0}(237,259)(216,259)(216,225){1}
wire [29:0] w0;    //: /sn:0 /dp:1 {0}(139,200)(191,200){1}
//: enddecls

  //: input g4 (WriteData) @(191,82) /sn:0 /w:[ 0 ]
  //: joint g8 (MemWrite) @(209, 124) /w:[ 2 1 -1 4 ]
  //: input g3 (MemWrite) @(149,111) /sn:0 /w:[ 0 ]
  tran g2(.Z(w0), .I(Address[31:2]));   //: @(133,200) /sn:0 /R:2 /w:[ 0 1 2 ] /ss:1
  //: input g1 (Address) @(86,213) /sn:0 /w:[ 0 ]
  //: comment g11 /dolink:0 /link:"" @(254,198) /sn:0
  //: /line:"D "
  //: /line:"(Read (1) de Lectura"
  //: /line:"(Write(1) de Escritura"
  //: /end
  //: supply0 g10 (w1) @(202,270) /sn:0 /w:[ 0 ]
  bufif1 g6 (.Z(ReadData), .I(WriteData), .E(MemWrite));   //: @(259,140) /sn:0 /w:[ 0 1 3 ]
  //: joint g7 (ReadData) @(277, 198) /w:[ 2 1 4 -1 ]
  //: input g9 (MemRead) @(239,259) /sn:0 /R:2 /w:[ 0 ]
  //: output g5 (ReadData) @(303,198) /sn:0 /w:[ 3 ]
  ram g0 (.A(w0), .D(ReadData), .WE(!MemWrite), .OE(!MemRead), .CS(w1));   //: @(209,199) /sn:0 /w:[ 1 5 5 1 1 ]
  //: comment g12 /dolink:0 /link:"" @(249,102) /sn:0
  //: /line:"Leer o Escribir"
  //: /end

endmodule

module SignExtend16to32bits(Adr32, Adr16);
//: interface  /sz:(156, 60) /bd:[ Ti0>Adr16[15:0](81/156) Ti1>Adr16[15:0](81/156) Bo0<Adr32[31:0](81/156) Bo1<Adr32[31:0](81/156) ]
input [15:0] Adr16;    //: /sn:0 {0}(220,171)(290,171){1}
//: {2}(291,171)(417,171){3}
supply1 [15:0] w43;    //: /sn:0 {0}(292,109)(292,145)(321,145){1}
output [31:0] Adr32;    //: /sn:0 /dp:1 {0}(423,166)(467,166){1}
wire [15:0] w45;    //: /sn:0 {0}(342,148)(353,148)(353,161)(417,161){1}
wire w39;    //: /sn:0 {0}(291,166)(291,150)(321,150){1}
//: enddecls

  //: supply1 g76 (w43) @(303,109) /sn:0 /w:[ 0 ]
  concat g72 (.I0(Adr16), .I1(w45), .Z(Adr32));   //: @(422,166) /sn:0 /w:[ 3 1 0 ] /dr:0
  //: output g1 (Adr32) @(464,166) /sn:0 /w:[ 1 ]
  tran g75(.Z(w39), .I(Adr16[15]));   //: @(291,169) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  and g74 (.I0(w43), .I1(w39), .Z(w45));   //: @(332,148) /sn:0 /w:[ 1 1 0 ]
  //: input g0 (Adr16) @(218,171) /sn:0 /w:[ 0 ]

endmodule

module Reg_16bits(D1, Clear, SelW, R1, Sel2, R2, D2, Wd, Clock, Wr, Sel1);
//: interface  /sz:(128, 88) /bd:[ Ti0>Clock(32/128) Ti1>Clear(107/128) Ti2>Clock(32/128) Ti3>Clear(107/128) Li0>SelW(83/88) Li1>Sel2(72/88) Li2>Sel1(60/88) Li3>Wr[3:0](46/88) Li4>R2[3:0](30/88) Li5>R1[3:0](16/88) Li6>SelW(83/88) Li7>Sel2(72/88) Li8>Sel1(60/88) Li9>Wr[3:0](46/88) Li10>R2[3:0](30/88) Li11>R1[3:0](16/88) Bi0>Wd[31:0](51/128) Bi1>Wd[31:0](51/128) Ri0>D2[31:0](60/88) Ri1>D1[31:0](20/88) Ri2>D2[31:0](60/88) Ri3>D1[31:0](20/88) ]
input [31:0] Wd;    //: /sn:0 /dp:1 {0}(339,387)(387,387){1}
//: {2}(391,387)(544,387){3}
//: {4}(548,387)(702,387){5}
//: {6}(706,387)(864,387)(864,363){7}
//: {8}(704,385)(704,267){9}
//: {10}(546,385)(546,154){11}
//: {12}(389,385)(389,39){13}
input Clock;    //: /sn:0 {0}(392,-82)(451,-82){1}
//: {2}(455,-82)(600,-82){3}
//: {4}(604,-82)(768,-82){5}
//: {6}(772,-82)(928,-82)(928,275){7}
//: {8}(770,-80)(770,179){9}
//: {10}(602,-80)(602,66){11}
//: {12}(453,-80)(453,-49){13}
output [31:0] D1;    //: /sn:0 /dp:1 {0}(952,303)(1077,303)(1077,204){1}
//: {2}(1077,200)(1077,87){3}
//: {4}(1077,83)(1077,-25){5}
//: {6}(1077,-29)(1077,-52)(1167,-52){7}
//: {8}(1075,-27)(476,-27){9}
//: {10}(1075,85)(629,85){11}
//: {12}(1075,202)(789,202){13}
output [31:0] D2;    //: /sn:0 /dp:13 {0}(952,338)(1120,338)(1120,252){1}
//: {2}(1120,248)(1120,132){3}
//: {4}(1120,128)(1120,18){5}
//: {6}(1120,14)(1120,-28)(1168,-28){7}
//: {8}(1118,16)(476,16){9}
//: {10}(1118,130)(629,130){11}
//: {12}(1118,250)(789,250){13}
input Clear;    //: /sn:0 {0}(393,-64)(399,-64){1}
//: {2}(403,-64)(541,-64){3}
//: {4}(545,-64)(697,-64){5}
//: {6}(701,-64)(868,-64)(868,275){7}
//: {8}(699,-62)(699,179){9}
//: {10}(543,-62)(543,66){11}
//: {12}(401,-62)(401,-49){13}
input [3:0] R2;    //: /sn:0 {0}(178,-69)(178,-17){1}
//: {2}(178,-16)(178,170){3}
//: {4}(178,171)(178,178){5}
input Sel2;    //: /sn:0 {0}(101,206)(244,206)(244,193){1}
input [3:0] Wr;    //: /sn:0 {0}(206,-70)(206,-2){1}
//: {2}(206,-1)(206,267){3}
//: {4}(206,268)(206,273){5}
input [3:0] R1;    //: /sn:0 {0}(150,-69)(150,-37){1}
//: {2}(150,-36)(150,60){3}
//: {4}(150,61)(150,66){5}
input SelW;    //: /sn:0 {0}(104,306)(249,306)(249,290){1}
input Sel1;    //: /sn:0 {0}(98,108)(238,108)(238,83){1}
wire w6;    //: /sn:0 {0}(254,67)(649,67)(649,237)(659,237){1}
wire w7;    //: /sn:0 {0}(254,55)(489,55)(489,128)(499,128){1}
wire w14;    //: /sn:0 {0}(260,153)(329,153)(329,20)(346,20){1}
wire [1:0] w15;    //: /sn:0 {0}(210,268)(236,268){1}
wire w19;    //: /sn:0 {0}(265,262)(484,262)(484,145)(499,145){1}
wire [1:0] w0;    //: /sn:0 {0}(154,-36)(309,-36){1}
//: {2}(313,-36)(346,-36){3}
//: {4}(311,-34)(311,82)(478,82){5}
//: {6}(482,82)(499,82){7}
//: {8}(480,84)(480,196)(627,196){9}
//: {10}(631,196)(659,196){11}
//: {12}(629,198)(629,288)(822,288){13}
wire [1:0] w3;    //: /sn:0 {0}(154,61)(225,61){1}
wire w20;    //: /sn:0 {0}(265,250)(322,250)(322,28)(346,28){1}
wire [1:0] w1;    //: /sn:0 {0}(182,-16)(295,-16){1}
//: {2}(299,-16)(346,-16){3}
//: {4}(297,-14)(297,97)(463,97){5}
//: {6}(467,97)(499,97){7}
//: {8}(465,99)(465,211)(613,211){9}
//: {10}(617,211)(659,211){11}
//: {12}(615,213)(615,305)(822,305){13}
wire w8;    //: /sn:0 {0}(254,43)(336,43)(336,11)(346,11){1}
wire w18;    //: /sn:0 {0}(265,274)(649,274)(649,258)(659,258){1}
wire w17;    //: /sn:0 {0}(265,286)(583,286)(583,356)(822,356){1}
wire [1:0] w22;    //: /sn:0 {0}(182,171)(231,171){1}
wire [1:0] w2;    //: /sn:0 /dp:1 {0}(210,-1)(282,-1){1}
//: {2}(286,-1)(346,-1){3}
//: {4}(284,1)(284,114)(453,114){5}
//: {6}(457,114)(499,114){7}
//: {8}(455,116)(455,223)(604,223){9}
//: {10}(608,223)(659,223){11}
//: {12}(606,225)(606,319)(822,319){13}
wire w11;    //: /sn:0 {0}(260,189)(628,189)(628,165)(809,165)(809,343)(822,343){1}
wire w12;    //: /sn:0 {0}(260,177)(641,177)(641,247)(659,247){1}
wire w13;    //: /sn:0 {0}(260,165)(489,165)(489,136)(499,136){1}
wire w5;    //: /sn:0 {0}(254,79)(497,79)(497,52)(801,52)(801,332)(822,332){1}
//: enddecls

  //: output g4 (D1) @(1164,-52) /sn:0 /w:[ 7 ]
  //: joint g8 (D1) @(1077, 202) /w:[ -1 2 12 1 ]
  Reg_4bits g3 (.CLR(Clear), .CLOCK(Clock), .SelW(w17), .Sel2(w11), .Sel1(w5), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(823, 276) /sz:(128, 86) /sn:0 /p:[ Ti0>7 Ti1>7 Li0>1 Li1>1 Li2>1 Li3>13 Li4>13 Li5>13 Bi0>7 Ro0<0 Ro1<0 ]
  //: input g13 (Clear) @(391,-64) /sn:0 /w:[ 0 ]
  //: joint g34 (w0) @(311, -36) /w:[ 2 -1 1 4 ]
  //: joint g37 (w1) @(297, -16) /w:[ 2 -1 1 4 ]
  //: input g51 (SelW) @(102,306) /sn:0 /w:[ 0 ]
  Reg_4bits g2 (.CLR(Clear), .CLOCK(Clock), .SelW(w18), .Sel2(w12), .Sel1(w6), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(660, 180) /sz:(128, 86) /sn:0 /p:[ Ti0>9 Ti1>9 Li0>1 Li1>1 Li2>1 Li3>11 Li4>11 Li5>11 Bi0>9 Ro0<13 Ro1<13 ]
  Reg_4bits g1 (.CLR(Clear), .CLOCK(Clock), .SelW(w19), .Sel2(w13), .Sel1(w7), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(500, 67) /sz:(128, 86) /sn:0 /p:[ Ti0>11 Ti1>11 Li0>1 Li1>1 Li2>1 Li3>7 Li4>7 Li5>7 Bi0>11 Ro0<11 Ro1<11 ]
  //: joint g11 (D2) @(1120, 16) /w:[ -1 6 8 5 ]
  //: joint g16 (Clock) @(453, -82) /w:[ 2 -1 1 12 ]
  //: joint g10 (D2) @(1120, 130) /w:[ -1 4 10 3 ]
  //: input g28 (R1) @(150,-71) /sn:0 /R:3 /w:[ 0 ]
  //: input g50 (Sel2) @(99,206) /sn:0 /w:[ 0 ]
  //: joint g19 (Clear) @(543, -64) /w:[ 4 -1 3 10 ]
  //: joint g27 (Wd) @(389, 387) /w:[ 2 12 1 -1 ]
  tran g32(.Z(w1), .I(R2[1:0]));   //: @(176,-16) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g6 (D1) @(1077, -27) /w:[ -1 6 8 5 ]
  //: joint g38 (w1) @(465, 97) /w:[ 6 -1 5 8 ]
  //: joint g7 (D1) @(1077, 85) /w:[ -1 4 10 3 ]
  //: joint g9 (D2) @(1120, 250) /w:[ -1 2 12 1 ]
  //: joint g15 (Clock) @(602, -82) /w:[ 4 -1 3 10 ]
  tran g31(.Z(w0), .I(R1[1:0]));   //: @(148,-36) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g39 (w1) @(615, 211) /w:[ 10 -1 9 12 ]
  demux g43 (.I(w3), .E(Sel1), .Z0(w5), .Z1(w6), .Z2(w7), .Z3(w8));   //: @(238,61) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 ]
  tran g48(.Z(w15), .I(Wr[3:2]));   //: @(204,268) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g17 (Clear) @(401, -64) /w:[ 2 -1 1 12 ]
  //: joint g25 (Wd) @(704, 387) /w:[ 6 8 5 -1 ]
  //: input g29 (R2) @(178,-71) /sn:0 /R:3 /w:[ 0 ]
  //: joint g42 (w2) @(606, 223) /w:[ 10 -1 9 12 ]
  //: output g5 (D2) @(1165,-28) /sn:0 /w:[ 7 ]
  //: joint g14 (Clock) @(770, -82) /w:[ 6 -1 5 8 ]
  tran g44(.Z(w3), .I(R1[3:2]));   //: @(148,61) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  demux g47 (.I(w15), .E(SelW), .Z0(w17), .Z1(w18), .Z2(w19), .Z3(w20));   //: @(249,268) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 ]
  //: input g24 (Wd) @(337,387) /sn:0 /w:[ 0 ]
  //: joint g36 (w0) @(629, 196) /w:[ 10 -1 9 12 ]
  //: joint g41 (w2) @(455, 114) /w:[ 6 -1 5 8 ]
  //: joint g40 (w2) @(284, -1) /w:[ 2 -1 1 4 ]
  Reg_4bits g0 (.CLOCK(Clock), .CLR(Clear), .SelW(w20), .Sel2(w14), .Sel1(w8), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(347, -48) /sz:(128, 86) /sn:0 /p:[ Ti0>13 Ti1>13 Li0>1 Li1>1 Li2>1 Li3>3 Li4>3 Li5>3 Bi0>13 Ro0<9 Ro1<9 ]
  //: joint g26 (Wd) @(546, 387) /w:[ 4 10 3 -1 ]
  //: joint g35 (w0) @(480, 82) /w:[ 6 -1 5 8 ]
  demux g45 (.I(w22), .E(Sel2), .Z0(w11), .Z1(w12), .Z2(w13), .Z3(w14));   //: @(244,171) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 ]
  tran g46(.Z(w22), .I(R2[3:2]));   //: @(176,171) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: input g12 (Clock) @(390,-82) /sn:0 /w:[ 0 ]
  //: joint g18 (Clear) @(699, -64) /w:[ 6 -1 5 8 ]
  //: input g30 (Wr) @(206,-72) /sn:0 /R:3 /w:[ 0 ]
  tran g33(.Z(w2), .I(Wr[1:0]));   //: @(204,-1) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g49 (Sel1) @(96,108) /sn:0 /w:[ 0 ]

endmodule

module Reg_32bits(R2, RegWrite, Wr, Clock, Clear, D1, D2, Wd, R1);
//: interface  /sz:(124, 113) /bd:[ Ti0>Clock(89/124) Ti1>Clear(38/124) Ti2>Clock(89/124) Ti3>Clear(38/124) Li0>R1[4:0](35/113) Li1>R2[4:0](49/113) Li2>Wr[4:0](18/113) Li3>R1[4:0](35/113) Li4>R2[4:0](49/113) Li5>Wr[4:0](18/113) Bi0>Wd[31:0](40/124) Bi1>RegWrite(92/124) Bi2>Wd[31:0](40/124) Bi3>RegWrite(92/124) Ro0<D2[31:0](73/113) Ro1<D1[31:0](41/113) Ro2<D2[31:0](73/113) Ro3<D1[31:0](41/113) ]
input [31:0] Wd;    //: /sn:0 /dp:1 {0}(639,192)(639,436)(522,436){1}
//: {2}(520,434)(520,399){3}
//: {4}(518,436)(375,436){5}
input Clock;    //: /sn:0 {0}(487,46)(557,46){1}
//: {2}(561,46)(620,46)(620,102){3}
//: {4}(559,48)(559,309){5}
supply1 w4;    //: /sn:0 {0}(177,322)(366,322)(366,312){1}
output [31:0] D1;    //: /sn:0 /dp:1 {0}(717,123)(829,123)(829,328){1}
//: {2}(827,330)(600,330){3}
//: {4}(829,332)(829,408)(868,408){5}
output [31:0] D2;    //: /sn:0 /dp:1 {0}(717,163)(779,163)(779,379){1}
//: {2}(777,381)(600,381){3}
//: {4}(779,383)(779,430)(868,430){5}
input Clear;    //: /sn:0 {0}(488,28)(514,28){1}
//: {2}(518,28)(695,28)(695,102){3}
//: {4}(516,30)(516,309){5}
input [4:0] R2;    //: /sn:0 {0}(292,102)(292,132){1}
//: {2}(292,133)(292,287){3}
//: {4}(292,288)(292,296){5}
input [4:0] Wr;    //: /sn:0 {0}(324,100)(324,149){1}
//: {2}(324,150)(324,361){3}
//: {4}(324,362)(324,367){5}
input [4:0] R1;    //: /sn:0 {0}(263,102)(263,118){1}
//: {2}(263,119)(263,200){3}
//: {4}(263,201)(263,207){5}
supply1 w12;    //: /sn:0 {0}(177,241)(363,241)(363,225){1}
input RegWrite;    //: /sn:0 {0}(229,409)(369,409)(369,385){1}
wire w6;    //: /sn:0 {0}(379,193)(540,193)(540,163)(587,163){1}
wire w7;    //: /sn:0 {0}(296,288)(304,288)(304,290)(353,290){1}
wire w14;    //: /sn:0 {0}(385,353)(421,353)(421,186)(587,186){1}
wire [3:0] w0;    //: /sn:0 {0}(267,119)(456,119){1}
//: {2}(460,119)(587,119){3}
//: {4}(458,121)(458,321)(470,321){5}
wire w3;    //: /sn:0 {0}(267,201)(275,201)(275,203)(350,203){1}
wire [3:0] w1;    //: /sn:0 {0}(296,133)(427,133){1}
//: {2}(431,133)(587,133){3}
//: {4}(429,135)(429,331)(470,331){5}
wire [3:0] w2;    //: /sn:0 {0}(328,150)(334,150)(334,149)(406,149){1}
//: {2}(410,149)(587,149){3}
//: {4}(408,151)(408,346)(470,346){5}
wire w11;    //: /sn:0 {0}(328,362)(336,362)(336,363)(356,363){1}
wire w10;    //: /sn:0 {0}(382,280)(550,280)(550,175)(587,175){1}
wire w13;    //: /sn:0 {0}(385,373)(450,373)(450,391)(470,391){1}
wire w5;    //: /sn:0 {0}(379,213)(449,213)(449,363)(470,363){1}
wire w9;    //: /sn:0 {0}(382,300)(460,300)(460,378)(470,378){1}
//: enddecls

  //: input g4 (R2) @(292,100) /sn:0 /R:3 /w:[ 0 ]
  //: input g8 (RegWrite) @(227,409) /sn:0 /w:[ 0 ]
  //: input g3 (Wr) @(324,98) /sn:0 /R:3 /w:[ 0 ]
  //: supply1 g13 (w12) @(177,230) /sn:0 /R:1 /w:[ 0 ]
  //: comment g34 /dolink:0 /link:"" @(920,398) /sn:0
  //: /line:"Salida, Contenido de los Reg's Selector's"
  //: /line:"R1 -> A (D1)"
  //: /line:"R2 -> B (D2)"
  //: /end
  //: joint g2 (Clear) @(516, 28) /w:[ 2 -1 1 4 ]
  Reg_16bits g1 (.Clock(Clock), .Clear(Clear), .SelW(w13), .Sel2(w9), .Sel1(w5), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(471, 310) /sz:(128, 88) /sn:0 /p:[ Ti0>5 Ti1>5 Li0>1 Li1>1 Li2>1 Li3>5 Li4>5 Li5>5 Bi0>3 Ri0>3 Ri1>3 ]
  //: input g11 (Clock) @(485,46) /sn:0 /w:[ 0 ]
  //: joint g16 (D2) @(779, 381) /w:[ -1 1 2 4 ]
  //: input g10 (Clear) @(486,28) /sn:0 /w:[ 0 ]
  tran g28(.Z(w11), .I(Wr[4]));   //: @(322,362) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g19(.Z(w1), .I(R2[3:0]));   //: @(290,133) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  tran g27(.Z(w7), .I(R2[4]));   //: @(290,288) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: comment g32 /dolink:0 /link:"" @(246,445) /sn:0
  //: /line:"Datos a Escribir al Reg a Modificar"
  //: /end
  //: output g6 (D1) @(865,408) /sn:0 /w:[ 5 ]
  //: output g7 (D2) @(865,430) /sn:0 /w:[ 5 ]
  //: input g9 (Wd) @(373,436) /sn:0 /w:[ 5 ]
  //: joint g15 (D1) @(829, 330) /w:[ -1 1 2 4 ]
  //: joint g20 (w1) @(429, 133) /w:[ 2 -1 1 4 ]
  //: comment g31 /dolink:0 /link:"" @(92,379) /sn:0
  //: /line:"Seleciona Reg a Modificar"
  //: /end
  tran g17(.Z(w0), .I(R1[3:0]));   //: @(261,119) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  demux g25 (.I(w11), .E(RegWrite), .Z0(w13), .Z1(w14));   //: @(369,363) /sn:0 /R:1 /w:[ 1 1 0 0 ]
  //: supply1 g29 (w4) @(177,311) /sn:0 /R:1 /w:[ 0 ]
  //: input g5 (R1) @(263,100) /sn:0 /R:3 /w:[ 0 ]
  //: joint g14 (Wd) @(520, 436) /w:[ 1 2 4 -1 ]
  tran g21(.Z(w2), .I(Wr[3:0]));   //: @(322,150) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  demux g24 (.I(w7), .E(w4), .Z0(w9), .Z1(w10));   //: @(366,290) /sn:0 /R:1 /w:[ 1 1 0 0 ]
  demux g23 (.I(w3), .E(w12), .Z0(w5), .Z1(w6));   //: @(363,203) /sn:0 /R:1 /w:[ 1 1 0 0 ]
  Reg_16bits g0 (.Clock(Clock), .Clear(Clear), .SelW(w14), .Sel2(w10), .Sel1(w6), .Wr(w2), .R2(w1), .R1(w0), .Wd(Wd), .D2(D2), .D1(D1));   //: @(588, 103) /sz:(128, 88) /sn:0 /p:[ Ti0>3 Ti1>3 Li0>1 Li1>1 Li2>1 Li3>3 Li4>3 Li5>3 Bi0>0 Ri0>0 Ri1>0 ]
  //: joint g22 (w2) @(408, 149) /w:[ 2 -1 1 4 ]
  tran g26(.Z(w3), .I(R1[4]));   //: @(261,201) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: joint g12 (Clock) @(559, 46) /w:[ 2 -1 1 4 ]
  //: joint g18 (w0) @(458, 119) /w:[ 2 -1 1 4 ]
  //: comment g30 /dolink:0 /link:"" @(93,269) /sn:0
  //: /line:"Seleciona Reg a Leer"
  //: /end
  //: comment g33 /dolink:0 /link:"" @(245,62) /sn:0
  //: /line:"Reg's Selector's"
  //: /end

endmodule

module ALU(Z, B, ALUop, R, A);
//: interface  /sz:(60, 101) /bd:[ Ti0>ALUop[2:0](27/60) Ti1>ALUop[2:0](27/60) Li0>B[31:0](66/101) Li1>A[31:0](27/101) Li2>B[31:0](66/101) Li3>A[31:0](27/101) Ro0<Z(35/101) Ro1<R[31:0](59/101) Ro2<Z(35/101) Ro3<R[31:0](59/101) ]
supply0 [31:0] w6;    //: /sn:0 /dp:1 {0}(586,227)(358,227)(358,224)(348,224){1}
//: {2}(344,224)(334,224)(334,263){3}
//: {4}(336,265)(341,265)(341,292){5}
//: {6}(334,267)(334,292){7}
//: {8}(346,226)(346,236)(348,236)(348,292){9}
input [31:0] B;    //: /sn:0 {0}(104,91)(234,91){1}
//: {2}(238,91)(308,91)(308,119){3}
//: {4}(310,121)(347,121)(347,174){5}
//: {6}(308,123)(308,141)(311,141)(311,162){7}
//: {8}(236,93)(236,112)(253,112){9}
input [2:0] ALUop;    //: /sn:0 {0}(259,308)(280,308){1}
//: {2}(281,308)(315,308){3}
input [31:0] A;    //: /sn:0 /dp:1 {0}(316,162)(316,127)(313,127)(313,94){1}
//: {2}(315,92)(352,92)(352,174){3}
//: {4}(313,90)(313,59)(202,59){5}
//: {6}(198,59)(105,59){7}
//: {8}(200,61)(200,71)(204,71)(204,188){9}
output Z;    //: /sn:0 /dp:1 {0}(244,412)(249,412)(249,452)(286,452){1}
output [31:0] R;    //: /sn:0 {0}(418,374)(338,374)(338,321){1}
supply0 [30:0] w8;    //: /sn:0 {0}(419,308)(419,270)(405,270){1}
wire w4;    //: /sn:0 {0}(164,202)(154,202){1}
wire [31:0] w19;    //: /sn:0 {0}(349,195)(349,205)(321,205)(321,292){1}
wire w3;    //: /sn:0 {0}(281,303)(281,202)(240,202){1}
//: {2}(238,200)(238,117)(253,117){3}
//: {4}(236,202)(212,202){5}
wire w1;    //: /sn:0 {0}(332,258)(340,258)(340,245)(415,245)(415,260)(405,260){1}
wire [31:0] w25;    //: /sn:0 {0}(274,115)(284,115)(284,130)(172,130)(172,188){1}
wire [31:0] w12;    //: /sn:0 /dp:1 {0}(361,292)(361,265)(399,265){1}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(223,412)(188,412)(188,277){1}
//: {2}(190,275)(354,275)(354,292){3}
//: {4}(188,273)(188,253){5}
//: {6}(190,251)(328,251)(328,257){7}
//: {8}(328,258)(328,292){9}
//: {10}(188,249)(188,217){11}
wire [31:0] w5;    //: /sn:0 /dp:1 {0}(314,292)(314,193)(313,193)(313,183){1}
//: enddecls

  //: output g4 (Z) @(283,452) /sn:0 /w:[ 1 ]
  xor g8 (.I0(B), .I1(w3), .Z(w25));   //: @(264,115) /sn:0 /w:[ 9 3 0 ]
  mux g3 (.I0(w5), .I1(w19), .I2(w2), .I3(w6), .I4(w6), .I5(w6), .I6(w2), .I7(w12), .S(ALUop), .Z(R));   //: @(338,308) /sn:0 /w:[ 0 1 9 7 5 9 3 0 3 1 ] /ss:0 /do:0
  //: joint g13 (A) @(313, 92) /w:[ 2 4 -1 1 ]
  add g2 (.A(w25), .B(A), .S(w2), .CI(w3), .CO(w4));   //: @(188,204) /sn:0 /w:[ 1 9 11 5 0 ]
  //: input g1 (B) @(102,91) /sn:0 /w:[ 0 ]
  //: input g11 (ALUop) @(257,308) /sn:0 /w:[ 0 ]
  tran g16(.Z(w3), .I(ALUop[2]));   //: @(281,306) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  //: output g10 (R) @(415,374) /sn:0 /w:[ 0 ]
  //: joint g19 (w3) @(238, 202) /w:[ 1 2 4 -1 ]
  or g6 (.I0(A), .I1(B), .Z(w19));   //: @(349,185) /sn:0 /R:3 /w:[ 3 5 0 ]
  and g7 (.I0(A), .I1(B), .Z(w5));   //: @(313,173) /sn:0 /R:3 /w:[ 0 7 1 ]
  //: joint g9 (w2) @(188, 251) /w:[ 6 10 -1 5 ]
  //: joint g15 (B) @(236, 91) /w:[ 2 -1 1 8 ]
  //: joint g17 (w6) @(334, 265) /w:[ 4 3 -1 6 ]
  //: supply0 g25 (w6) @(592,227) /sn:0 /R:1 /w:[ 0 ]
  nor g5 (.I0(w2), .Z(Z));   //: @(234,412) /sn:0 /w:[ 0 0 ]
  //: joint g14 (A) @(200, 59) /w:[ 5 -1 6 8 ]
  concat g21 (.I0(w1), .I1(w8), .Z(w12));   //: @(400,265) /sn:0 /R:2 /w:[ 1 1 1 ] /dr:0
  //: joint g24 (w2) @(188, 275) /w:[ 2 4 -1 1 ]
  tran g23(.Z(w1), .I(w2[31]));   //: @(326,258) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: input g0 (A) @(103,59) /sn:0 /w:[ 7 ]
  //: supply0 g26 (w8) @(419,314) /sn:0 /w:[ 0 ]
  //: joint g12 (B) @(308, 121) /w:[ 4 3 -1 6 ]
  //: joint g18 (w6) @(346, 224) /w:[ 1 -1 2 8 ]

endmodule

module CONTROL(op, Branch, MemToReg, ALUsrc, MemRead, RegWrite, ALUop, Jump, MemWrite, RegDst);
//: interface  /sz:(941, 41) /bd:[ Bi0>op[5:0](870/941) Bi1>op[5:0](408/941) Bo0<Jump(710/941) Bo1<Branch(88/941) Bo2<RegDst(151/941) Bo3<ALUsrc(300/941) Bo4<RegWrite(220/941) Bo5<ALUop[1:0](370/941) Bo6<MemRead(620/941) Bo7<MemWrite(460/941) Bo8<MemToReg(530/941) ]
output MemToReg;    //: /sn:0 /dp:1 {0}(295,436)(354,436)(354,437)(693,437){1}
output [1:0] ALUop;    //: /sn:0 {0}(656,481)(700,481){1}
output Jump;    //: /sn:0 /dp:1 {0}(491,342)(491,627)(703,627){1}
output MemWrite;    //: /sn:0 /dp:1 {0}(305,343)(305,514){1}
//: {2}(307,516)(317,516)(317,517)(697,517){3}
//: {4}(305,518)(305,551){5}
//: {6}(307,553)(331,553)(331,540)(698,540){7}
//: {8}(305,555)(305,638){9}
output Branch;    //: /sn:0 /dp:1 {0}(396,630)(396,487){1}
//: {2}(398,485)(408,485)(408,486)(650,486){3}
//: {4}(396,483)(396,394){5}
//: {6}(398,392)(693,392){7}
//: {8}(396,390)(396,344){9}
output ALUsrc;    //: /sn:0 {0}(719,538)(737,538)(737,540)(846,540){1}
output RegDst;    //: /sn:0 {0}(694,582)(132,582){1}
//: {2}(130,580)(130,477){3}
//: {4}(132,475)(142,475)(142,476)(650,476){5}
//: {6}(130,473)(130,378){7}
//: {8}(132,376)(694,376){9}
//: {10}(130,374)(130,341){11}
//: {12}(130,584)(130,679){13}
output RegWrite;    //: /sn:0 /dp:1 {0}(715,585)(768,585)(768,581)(847,581){1}
input [5:0] op;    //: /sn:0 {0}(22,25)(50,25)(50,34){1}
//: {2}(50,35)(50,50){3}
//: {4}(50,51)(50,64){5}
//: {6}(50,65)(50,77){7}
//: {8}(50,78)(50,90){9}
//: {10}(50,91)(50,106){11}
//: {12}(50,107)(50,120){13}
output MemRead;    //: /sn:0 /dp:1 {0}(218,645)(218,587){1}
//: {2}(220,585)(230,585)(230,587)(694,587){3}
//: {4}(218,583)(218,539){5}
//: {6}(220,537)(232,537)(232,535)(698,535){7}
//: {8}(218,535)(218,437){9}
//: {10}(220,435)(273,435)(273,436)(279,436){11}
//: {12}(218,433)(218,421){13}
//: {14}(220,419)(230,419)(230,421)(694,421){15}
//: {16}(218,417)(218,344){17}
wire w32;    //: /sn:0 {0}(393,259)(393,323){1}
wire w7;    //: /sn:0 {0}(488,321)(488,275){1}
wire w16;    //: /sn:0 {0}(131,238)(131,278)(132,278)(132,320){1}
wire w4;    //: /sn:0 {0}(122,261)(122,320){1}
wire w19;    //: /sn:0 {0}(297,270)(297,322){1}
wire w0;    //: /sn:0 {0}(54,107)(104,107){1}
//: {2}(108,107)(227,107){3}
//: {4}(231,107)(319,107){5}
//: {6}(323,107)(404,107){7}
//: {8}(408,107)(478,107)(478,321){9}
//: {10}(406,109)(406,119)(408,119)(408,286){11}
//: {12}(321,109)(321,119)(317,119)(317,322){13}
//: {14}(229,109)(229,119)(230,119)(230,323){15}
//: {16}(106,109)(106,119)(115,119)(115,265){17}
wire w34;    //: /sn:0 {0}(383,221)(383,323){1}
wire w21;    //: /sn:0 {0}(215,289)(215,323){1}
wire w31;    //: /sn:0 {0}(408,302)(408,323){1}
wire w28;    //: /sn:0 {0}(54,51)(132,51){1}
//: {2}(136,51)(220,51){3}
//: {4}(224,51)(298,51){5}
//: {6}(302,51)(378,51){7}
//: {8}(382,51)(498,51)(498,262){9}
//: {10}(380,53)(380,63)(388,63)(388,220){11}
//: {12}(300,53)(300,63)(297,63)(297,254){13}
//: {14}(222,53)(222,63)(210,63)(210,238){15}
//: {16}(134,53)(134,63)(136,63)(136,169){17}
wire w24;    //: /sn:0 {0}(54,78)(120,78){1}
//: {2}(124,78)(219,78){3}
//: {4}(223,78)(308,78){5}
//: {6}(312,78)(394,78){7}
//: {8}(398,78)(488,78)(488,259){9}
//: {10}(396,80)(396,90)(398,90)(398,323){11}
//: {12}(310,80)(310,90)(307,90)(307,282){13}
//: {14}(221,80)(221,90)(220,90)(220,294){15}
//: {16}(122,80)(122,90)(126,90)(126,208){17}
wire w20;    //: /sn:0 {0}(498,278)(498,321){1}
wire w36;    //: /sn:0 {0}(142,169)(142,320){1}
wire w23;    //: /sn:0 {0}(210,254)(210,323){1}
wire w1;    //: /sn:0 {0}(115,281)(115,310)(117,310)(117,320){1}
wire w25;    //: /sn:0 {0}(54,65)(125,65){1}
//: {2}(129,65)(207,65){3}
//: {4}(211,65)(305,65){5}
//: {6}(309,65)(387,65){7}
//: {8}(391,65)(493,65)(493,215){9}
//: {10}(389,67)(389,77)(393,77)(393,243){11}
//: {12}(307,67)(307,77)(302,77)(302,322){13}
//: {14}(209,67)(209,77)(215,77)(215,273){15}
//: {16}(127,67)(127,77)(131,77)(131,222){17}
wire w35;    //: /sn:0 /dp:1 {0}(503,321)(503,197){1}
wire w8;    //: /sn:0 {0}(483,321)(483,294){1}
wire w30;    //: /sn:0 /dp:1 {0}(54,35)(142,35){1}
//: {2}(146,35)(205,35){3}
//: {4}(209,35)(292,35){5}
//: {6}(296,35)(371,35){7}
//: {8}(375,35)(503,35)(503,181){9}
//: {10}(373,37)(373,47)(383,47)(383,205){11}
//: {12}(294,37)(294,47)(292,47)(292,322){13}
//: {14}(207,37)(207,47)(205,47)(205,323){15}
//: {16}(144,37)(144,47)(142,47)(142,153){17}
wire w22;    //: /sn:0 {0}(54,91)(112,91){1}
//: {2}(116,91)(226,91){3}
//: {4}(230,91)(315,91){5}
//: {6}(319,91)(401,91){7}
//: {8}(405,91)(483,91)(483,278){9}
//: {10}(403,93)(403,263){11}
//: {12}(317,93)(317,103)(312,103)(312,322){13}
//: {14}(228,93)(228,103)(225,103)(225,323){15}
//: {16}(114,93)(114,103)(122,103)(122,245){17}
wire w17;    //: /sn:0 {0}(493,231)(493,321){1}
wire w10;    //: /sn:0 {0}(126,224)(126,271)(127,271)(127,320){1}
wire w27;    //: /sn:0 {0}(136,185)(136,252)(137,252)(137,320){1}
wire w33;    //: /sn:0 {0}(388,236)(388,323){1}
wire w29;    //: /sn:0 {0}(403,279)(403,323){1}
wire w9;    //: /sn:0 {0}(307,298)(307,322){1}
wire w26;    //: /sn:0 {0}(220,310)(220,323){1}
//: enddecls

  tran g8(.Z(w28), .I(op[4]));   //: @(48,51) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: input g4 (op) @(20,25) /sn:0 /w:[ 0 ]
  //: joint g61 (MemRead) @(218, 435) /w:[ 10 12 -1 9 ]
  //: joint g58 (RegDst) @(130, 376) /w:[ 8 10 -1 7 ]
  //: output g55 (Branch) @(690,392) /sn:0 /w:[ 7 ]
  //: output g51 (MemToReg) @(690,437) /sn:0 /w:[ 1 ]
  not g37 (.I(w30), .Z(w36));   //: @(142,159) /sn:0 /R:3 /w:[ 17 0 ]
  not g34 (.I(w24), .Z(w10));   //: @(126,214) /sn:0 /R:3 /w:[ 17 0 ]
  tran g13(.Z(w22), .I(op[1]));   //: @(48,91) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  and g3 (.I0(w31), .I1(w29), .I2(w24), .I3(w32), .I4(w33), .I5(w34), .Z(Branch));   //: @(396,334) /sn:0 /R:3 /w:[ 1 1 11 1 1 1 9 ]
  //: joint g65 (RegDst) @(130, 475) /w:[ 4 6 -1 3 ]
  //: joint g77 (w28) @(222, 51) /w:[ 4 -1 3 14 ]
  //: joint g76 (w25) @(209, 65) /w:[ 4 -1 3 14 ]
  and g2 (.I0(w0), .I1(w22), .I2(w9), .I3(w25), .I4(w19), .I5(w30), .Z(MemWrite));   //: @(305,333) /sn:0 /R:3 /w:[ 13 13 1 13 1 13 0 ]
  //: joint g59 (Branch) @(396, 485) /w:[ 2 4 -1 1 ]
  and g72 (.I0(w35), .I1(w20), .I2(w17), .I3(w7), .I4(w8), .I5(w0), .Z(Jump));   //: @(491,332) /sn:0 /R:3 /w:[ 0 1 1 0 0 9 0 ]
  and g1 (.I0(w0), .I1(w22), .I2(w26), .I3(w21), .I4(w23), .I5(w30), .Z(MemRead));   //: @(218,334) /sn:0 /R:3 /w:[ 15 15 1 1 1 15 17 ]
  //: joint g64 (Branch) @(396, 392) /w:[ 6 8 -1 5 ]
  //: joint g16 (w0) @(406, 107) /w:[ 8 -1 7 10 ]
  tran g11(.Z(w24), .I(op[2]));   //: @(48,78) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: joint g78 (w30) @(207, 35) /w:[ 4 -1 3 14 ]
  //: joint g28 (w22) @(317, 91) /w:[ 6 -1 5 12 ]
  //: output g50 (ALUsrc) @(843,540) /sn:0 /w:[ 1 ]
  not g10 (.I(w25), .Z(w32));   //: @(393,249) /sn:0 /R:3 /w:[ 11 0 ]
  //: joint g32 (w30) @(294, 35) /w:[ 6 -1 5 12 ]
  //: joint g27 (w0) @(321, 107) /w:[ 6 -1 5 12 ]
  //: joint g19 (w24) @(396, 78) /w:[ 8 -1 7 10 ]
  //: joint g69 (RegDst) @(130, 582) /w:[ 1 2 -1 12 ]
  not g38 (.I(w0), .Z(w1));   //: @(115,271) /sn:0 /R:3 /w:[ 17 0 ]
  not g6 (.I(w0), .Z(w31));   //: @(408,292) /sn:0 /R:3 /w:[ 11 0 ]
  //: joint g75 (w24) @(221, 78) /w:[ 4 -1 3 14 ]
  concat g57 (.I0(Branch), .I1(RegDst), .Z(ALUop));   //: @(655,481) /sn:0 /w:[ 3 5 0 ] /dr:0
  //: output g53 (MemRead) @(691,421) /sn:0 /w:[ 15 ]
  tran g9(.Z(w25), .I(op[3]));   //: @(48,65) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  not g7 (.I(w22), .Z(w29));   //: @(403,269) /sn:0 /R:3 /w:[ 11 0 ]
  //: joint g31 (w28) @(300, 51) /w:[ 6 -1 5 12 ]
  //: joint g20 (w25) @(389, 65) /w:[ 8 -1 7 10 ]
  buf g71 (.I(MemRead), .Z(MemToReg));   //: @(285,436) /sn:0 /w:[ 11 0 ]
  tran g15(.Z(w0), .I(op[0]));   //: @(48,107) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  //: joint g68 (MemWrite) @(305, 553) /w:[ 6 5 -1 8 ]
  //: joint g67 (MemRead) @(218, 537) /w:[ 6 8 -1 5 ]
  //: joint g39 (w30) @(144, 35) /w:[ 2 -1 1 16 ]
  //: comment g48 /dolink:0 /link:"" @(363,339) /sn:0 /R:3
  //: /line:"BEQ"
  //: /end
  //: joint g43 (w22) @(114, 91) /w:[ 2 -1 1 16 ]
  //: joint g73 (w0) @(229, 107) /w:[ 4 -1 3 14 ]
  //: joint g29 (w24) @(310, 78) /w:[ 6 -1 5 12 ]
  //: joint g17 (w22) @(403, 91) /w:[ 8 -1 7 10 ]
  //: joint g62 (MemWrite) @(305, 516) /w:[ 2 1 -1 4 ]
  not g25 (.I(w28), .Z(w23));   //: @(210,244) /sn:0 /R:3 /w:[ 15 0 ]
  or g63 (.I0(RegDst), .I1(MemRead), .Z(RegWrite));   //: @(705,585) /sn:0 /w:[ 0 3 0 ]
  //: output g52 (RegWrite) @(844,581) /sn:0 /w:[ 1 ]
  //: joint g42 (w24) @(122, 78) /w:[ 2 -1 1 16 ]
  not g83 (.I(w24), .Z(w7));   //: @(488,265) /sn:0 /R:3 /w:[ 9 1 ]
  //: joint g74 (w22) @(228, 91) /w:[ 4 -1 3 14 ]
  //: output g56 (ALUop) @(697,481) /sn:0 /w:[ 1 ]
  not g14 (.I(w30), .Z(w34));   //: @(383,211) /sn:0 /R:3 /w:[ 11 0 ]
  tran g5(.Z(w30), .I(op[5]));   //: @(48,35) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: output g80 (Jump) @(700,627) /sn:0 /w:[ 1 ]
  //: comment g79 /dolink:0 /link:"" @(456,343) /sn:0
  //: /line:"Jump"
  //: /end
  //: comment g47 /dolink:0 /link:"" @(278,338) /sn:0 /R:3
  //: /line:"SW"
  //: /end
  //: joint g44 (w0) @(106, 107) /w:[ 2 -1 1 16 ]
  //: joint g24 (w30) @(373, 35) /w:[ 8 -1 7 10 ]
  not g85 (.I(w28), .Z(w20));   //: @(498,268) /sn:0 /R:3 /w:[ 9 0 ]
  not g84 (.I(w25), .Z(w17));   //: @(493,221) /sn:0 /R:3 /w:[ 9 0 ]
  not g36 (.I(w28), .Z(w27));   //: @(136,175) /sn:0 /R:3 /w:[ 17 0 ]
  not g21 (.I(w28), .Z(w19));   //: @(297,260) /sn:0 /R:3 /w:[ 13 0 ]
  //: joint g41 (w25) @(127, 65) /w:[ 2 -1 1 16 ]
  not g23 (.I(w25), .Z(w21));   //: @(215,279) /sn:0 /R:3 /w:[ 15 0 ]
  not g81 (.I(w22), .Z(w8));   //: @(483,284) /sn:0 /R:3 /w:[ 9 1 ]
  //: joint g60 (MemRead) @(218, 419) /w:[ 14 16 -1 13 ]
  //: output g54 (MemWrite) @(694,517) /sn:0 /w:[ 3 ]
  //: joint g40 (w28) @(134, 51) /w:[ 2 -1 1 16 ]
  //: joint g22 (w28) @(380, 51) /w:[ 8 -1 7 10 ]
  //: joint g70 (MemRead) @(218, 585) /w:[ 2 4 -1 1 ]
  //: comment g46 /dolink:0 /link:"" @(184,334) /sn:0 /R:3
  //: /line:"LW"
  //: /end
  //: comment g45 /dolink:0 /link:"" @(58,332) /sn:0 /R:3
  //: /line:"R-format"
  //: /end
  not g35 (.I(w25), .Z(w16));   //: @(131,228) /sn:0 /R:3 /w:[ 17 0 ]
  not g26 (.I(w24), .Z(w26));   //: @(220,300) /sn:0 /R:3 /w:[ 15 0 ]
  and g0 (.I0(w36), .I1(w27), .I2(w16), .I3(w10), .I4(w4), .I5(w1), .Z(RegDst));   //: @(130,331) /sn:0 /R:3 /w:[ 1 1 1 1 1 1 11 ]
  not g82 (.I(w30), .Z(w35));   //: @(503,187) /sn:0 /R:3 /w:[ 9 1 ]
  or g66 (.I0(MemRead), .I1(MemWrite), .Z(ALUsrc));   //: @(709,538) /sn:0 /w:[ 7 7 0 ]
  not g18 (.I(w24), .Z(w9));   //: @(307,288) /sn:0 /R:3 /w:[ 13 0 ]
  not g12 (.I(w28), .Z(w33));   //: @(388,226) /sn:0 /R:3 /w:[ 11 0 ]
  //: joint g30 (w25) @(307, 65) /w:[ 6 -1 5 12 ]
  not g33 (.I(w22), .Z(w4));   //: @(122,251) /sn:0 /R:3 /w:[ 17 0 ]
  //: output g49 (RegDst) @(691,376) /sn:0 /w:[ 9 ]

endmodule

module BEQ(Sum, Btarget, PC);
//: interface  /sz:(81, 100) /bd:[ Li0>PC[31:0](27/100) Li1>Btarget[31:0](75/100) Ro0<Sum[31:0](48/100) ]
input [31:0] Btarget;    //: /sn:0 {0}(144,187)(228,187)(228,304)(371,304)(371,269)(432,269)(432,196)(468,196){1}
input [31:0] PC;    //: /sn:0 {0}(314,151)(428,151)(428,164)(468,164){1}
supply0 w1;    //: /sn:0 {0}(482,127)(482,156){1}
output [31:0] Sum;    //: /sn:0 /dp:1 {0}(497,180)(598,180)(598,300)(629,300){1}
wire w6;    //: /sn:0 {0}(482,204)(482,214){1}
//: enddecls

  //: output g2 (Sum) @(626,300) /sn:0 /w:[ 1 ]
  //: input g1 (Btarget) @(142,187) /sn:0 /w:[ 0 ]
  add g6 (.A(Btarget), .B(PC), .S(Sum), .CI(w1), .CO(w6));   //: @(484,180) /sn:0 /R:1 /w:[ 1 1 0 1 0 ]
  //: supply0 g7 (w1) @(482,121) /sn:0 /R:2 /w:[ 0 ]
  //: input g0 (PC) @(312,151) /sn:0 /w:[ 0 ]

endmodule

module Reg_4bits(CLR, Sel1, R1, D2, D1, Wd, Wr, CLOCK, Sel2, SelW, R2);
//: interface  /sz:(128, 86) /bd:[ Ti0>CLR(39/128) Ti1>CLOCK(110/128) Ti2>CLR(39/128) Ti3>CLOCK(110/128) Li0>SelW(78/86) Li1>Sel2(67/86) Li2>Sel1(57/86) Li3>Wr[1:0](43/86) Li4>R2[1:0](31/86) Li5>R1[1:0](16/86) Li6>SelW(78/86) Li7>Sel2(67/86) Li8>Sel1(57/86) Li9>Wr[1:0](43/86) Li10>R2[1:0](31/86) Li11>R1[1:0](16/86) Bi0>Wd[31:0](44/128) Bi1>Wd[31:0](44/128) Ro0<D2[31:0](70/86) Ro1<D1[31:0](22/86) Ro2<D2[31:0](70/86) Ro3<D1[31:0](22/86) ]
input [31:0] Wd;    //: /sn:0 {0}(35,174)(144,174){1}
//: {2}(148,174)(237,174){3}
//: {4}(241,174)(340,174){5}
//: {6}(344,174)(443,174)(443,295){7}
//: {8}(342,176)(342,257){9}
//: {10}(239,176)(239,204)(239,204)(239,228){11}
//: {12}(146,176)(146,194){13}
output [31:0] D1;    //: /sn:0 {0}(422,467)(438,467)(438,497)(464,497){1}
output [31:0] D2;    //: /sn:0 {0}(281,498)(291,498)(291,522)(462,522){1}
input [1:0] R2;    //: /sn:0 /dp:1 {0}(-12,443)(188,443){1}
input Sel2;    //: /sn:0 {0}(263,466)(273,466)(273,493){1}
input [1:0] Wr;    //: /sn:0 {0}(553,166)(553,135)(33,135){1}
input CLR;    //: /sn:0 {0}(497,36)(497,197){1}
//: {2}(495,199)(185,199){3}
//: {4}(497,201)(497,231){5}
//: {6}(495,233)(278,233){7}
//: {8}(497,235)(497,260){9}
//: {10}(495,262)(381,262){11}
//: {12}(497,264)(497,300)(482,300){13}
input [1:0] R1;    //: /sn:0 {0}(-11,399)(317,399){1}
input SelW;    //: /sn:0 /dp:1 {0}(529,179)(518,179)(518,106)(449,106){1}
input Sel1;    //: /sn:0 {0}(398,437)(414,437)(414,462){1}
input CLOCK;    //: /sn:0 {0}(-32,52)(-32,202){1}
//: {2}(-30,204)(109,204){3}
//: {4}(-32,206)(-32,236){5}
//: {6}(-30,238)(202,238){7}
//: {8}(-32,240)(-32,265){9}
//: {10}(-30,267)(305,267){11}
//: {12}(-32,269)(-32,305)(406,305){13}
wire [31:0] w15;    //: /sn:0 {0}(443,316)(443,346)(351,346)(351,367){1}
//: {2}(353,369)(358,369)(358,383){3}
//: {4}(349,369)(229,369)(229,427){5}
wire [31:0] w0;    //: /sn:0 {0}(146,215)(146,336)(219,336)(219,344){1}
//: {2}(221,346)(322,346)(322,383){3}
//: {4}(217,346)(193,346)(193,427){5}
wire w28;    //: /sn:0 {0}(559,195)(559,272)(381,272){1}
wire [31:0] w1;    //: /sn:0 {0}(340,412)(340,467)(406,467){1}
wire [31:0] w2;    //: /sn:0 {0}(211,456)(211,498)(265,498){1}
wire [31:0] w10;    //: /sn:0 {0}(342,278)(342,358){1}
//: {2}(344,360)(346,360)(346,383){3}
//: {4}(340,360)(217,360)(217,427){5}
wire w27;    //: /sn:0 {0}(547,195)(547,243)(278,243){1}
wire [31:0] w5;    //: /sn:0 {0}(239,249)(239,351){1}
//: {2}(241,353)(334,353)(334,383){3}
//: {4}(237,353)(205,353)(205,427){5}
wire w29;    //: /sn:0 {0}(571,195)(571,310)(482,310){1}
wire w26;    //: /sn:0 {0}(535,195)(535,209)(185,209){1}
//: enddecls

  mux g8 (.I0(w0), .I1(w5), .I2(w10), .I3(w15), .S(R2), .Z(w2));   //: @(211,443) /sn:0 /w:[ 5 5 5 5 1 0 ] /ss:0 /do:0
  //: input g4 (CLR) @(497,34) /sn:0 /R:3 /w:[ 0 ]
  register g3 (.Q(w15), .D(Wd), .EN(!w29), .CLR(!CLR), .CK(CLOCK));   //: @(443,305) /sn:0 /w:[ 0 7 1 13 13 ]
  //: joint g13 (w0) @(219, 346) /w:[ 2 1 4 -1 ]
  bufif1 g34 (.Z(D2), .I(w2), .E(Sel2));   //: @(271,498) /sn:0 /w:[ 0 1 1 ]
  //: input g37 (Sel1) @(396,437) /sn:0 /w:[ 0 ]
  register g2 (.Q(w10), .D(Wd), .EN(!w28), .CLR(!CLR), .CK(CLOCK));   //: @(342,267) /sn:0 /w:[ 0 9 1 11 11 ]
  register g1 (.Q(w5), .D(Wd), .EN(!w27), .CLR(!CLR), .CK(CLOCK));   //: @(239,238) /sn:0 /w:[ 0 11 1 7 7 ]
  //: input g11 (R1) @(-13,399) /sn:0 /w:[ 0 ]
  //: joint g16 (w15) @(351, 369) /w:[ 2 1 4 -1 ]
  mux g10 (.I0(w0), .I1(w5), .I2(w10), .I3(w15), .S(R1), .Z(w1));   //: @(340,399) /sn:0 /w:[ 3 3 3 3 1 0 ] /ss:0 /do:0
  //: output g28 (D2) @(459,522) /sn:0 /w:[ 1 ]
  //: joint g19 (Wd) @(342, 174) /w:[ 6 -1 5 8 ]
  //: output g27 (D1) @(461,497) /sn:0 /w:[ 1 ]
  //: comment g32 /dolink:0 /link:"" @(-109,412) /sn:0
  //: /line:"Registres a Seleccionar"
  //: /end
  //: joint g6 (CLR) @(497, 233) /w:[ -1 5 6 8 ]
  demux g9 (.I(Wr), .E(SelW), .Z0(w26), .Z1(w27), .Z2(w28), .Z3(w29));   //: @(553,179) /sn:0 /w:[ 0 0 0 0 0 0 ]
  //: joint g7 (CLR) @(497, 199) /w:[ -1 1 2 4 ]
  //: joint g15 (w10) @(342, 360) /w:[ 2 1 4 -1 ]
  //: joint g20 (Wd) @(146, 174) /w:[ 2 -1 1 12 ]
  //: comment g31 /dolink:0 /link:"" @(-22,145) /sn:0
  //: /line:"Dades a ficar al Registre"
  //: /end
  //: input g17 (Wd) @(33,174) /sn:0 /w:[ 0 ]
  //: input g25 (Wr) @(31,135) /sn:0 /w:[ 1 ]
  //: comment g29 /dolink:0 /link:"" @(389,86) /sn:0
  //: /line:"Control"
  //: /end
  //: joint g14 (w5) @(239, 353) /w:[ 2 1 4 -1 ]
  //: joint g5 (CLR) @(497, 262) /w:[ -1 9 10 12 ]
  //: input g21 (CLOCK) @(-32,50) /sn:0 /R:3 /w:[ 0 ]
  //: joint g24 (CLOCK) @(-32, 204) /w:[ 2 1 -1 4 ]
  //: input g36 (Sel2) @(261,466) /sn:0 /w:[ 0 ]
  //: joint g23 (CLOCK) @(-32, 238) /w:[ 6 5 -1 8 ]
  register g0 (.Q(w0), .D(Wd), .EN(!w26), .CLR(!CLR), .CK(CLOCK));   //: @(146,204) /sn:0 /w:[ 0 13 1 3 3 ]
  //: joint g22 (CLOCK) @(-32, 267) /w:[ 10 9 -1 12 ]
  //: input g26 (SelW) @(447,106) /sn:0 /w:[ 1 ]
  bufif1 g35 (.Z(D1), .I(w1), .E(Sel1));   //: @(412,467) /sn:0 /w:[ 0 1 1 ]
  //: input g12 (R2) @(-14,443) /sn:0 /w:[ 0 ]
  //: joint g18 (Wd) @(239, 174) /w:[ 4 -1 3 10 ]
  //: comment g30 /dolink:0 /link:"" @(-23,112) /sn:0
  //: /line:"Registre a Modificar"
  //: /end
  //: comment g33 /dolink:0 /link:"" @(384,501) /sn:0
  //: /line:"Dades Selecionats Sortida"
  //: /end

endmodule

module main;    //: root_module
supply0 w4;    //: /sn:0 {0}(-1149,523)(-1149,519)(-1249,519)(-1249,482){1}
supply0 w3;    //: /sn:0 {0}(-1170,333)(-1170,354){1}
supply0 w36;    //: /sn:0 /dp:1 {0}(635,470)(635,440)(640,440)(640,431){1}
supply0 w11;    //: /sn:0 /dp:1 {0}(-1340,409)(-1340,382)(-1348,382){1}
wire w6;    //: /sn:0 {0}(-976,23)(-976,43)(-1001,43){1}
//: {2}(-1003,41)(-1003,-12){3}
//: {4}(-1003,45)(-1003,239)(-1089,239){5}
wire w32;    //: /sn:0 {0}(-982,373)(-926,373)(-926,47){1}
//: {2}(-928,45)(-928,45){3}
//: {4}(-926,43)(-926,-12){5}
//: {6}(-924,45)(-905,45)(-905,24){7}
wire [31:0] w7;    //: /sn:0 {0}(-1155,378)(-1140,378){1}
//: {2}(-1139,378)(-1099,378){3}
//: {4}(-1095,378)(-1079,378)(-1079,345){5}
//: {6}(-1097,376)(-1097,157)(94,157)(94,237)(105,237){7}
wire w45;    //: /sn:0 {0}(628,281)(642,281)(642,328){1}
//: {2}(644,330)(694,330)(694,341){3}
//: {4}(642,332)(642,354)(647,354)(647,367){5}
//: {6}(649,369)(674,369)(674,358){7}
//: {8}(647,371)(647,381){9}
wire [4:0] w46;    //: /sn:0 /dp:1 {0}(-344,456)(-364,456){1}
wire [4:0] w14;    //: /sn:0 {0}(-724,450)(-724,396){1}
//: {2}(-722,394)(-648,394){3}
//: {4}(-724,392)(-724,217){5}
wire [5:0] w15;    //: /sn:0 {0}(-686,450)(-686,428){1}
//: {2}(-684,426)(-663,426){3}
//: {4}(-662,426)(-655,426)(-655,360)(-110,360){5}
//: {6}(-686,424)(-686,217){7}
wire w19;    //: /sn:0 /dp:1 {0}(-982,378)(-973,378)(-973,679)(227,679)(227,611){1}
wire w38;    //: /sn:0 /dp:1 {0}(790,17)(790,40)(830,40){1}
//: {2}(832,38)(832,-12){3}
//: {4}(832,42)(832,381)(765,381)(765,469)(750,469)(750,459){5}
wire [29:0] w0;    //: /sn:0 /dp:1 {0}(-1277,565)(-1289,565)(-1289,461){1}
wire [31:0] w37;    //: /sn:0 {0}(-507,656)(-507,671)(-319,671){1}
//: {2}(-315,671)(-76,671)(-76,567){3}
//: {4}(-74,565)(-50,565){5}
//: {6}(-76,563)(-76,285)(105,285){7}
//: {8}(-317,673)(-317,690){9}
wire w34;    //: /sn:0 /dp:1 {0}(-1066,329)(-1037,329)(-1037,375)(-1003,375){1}
wire [31:0] w43;    //: /sn:0 /dp:1 {0}(188,258)(202,258)(202,227)(234,227){1}
//: {2}(236,225)(236,139)(-1154,139)(-1154,353)(-1099,353)(-1099,345){3}
//: {4}(236,229)(236,298){5}
wire w21;    //: /sn:0 {0}(607,283)(570,283)(570,37){1}
//: {2}(570,33)(570,-12){3}
//: {4}(568,35)(547,35)(547,14){5}
wire w31;    //: /sn:0 /dp:1 {0}(-305,365)(-305,322)(67,322)(67,60)(-806,60){1}
//: {2}(-810,60)(-1324,60)(-1324,372)(-1348,372){3}
//: {4}(-808,62)(-808,170)(312,170)(312,158){5}
wire w28;    //: /sn:0 {0}(-34,598)(-34,613)(36,613)(36,33){1}
//: {2}(36,29)(36,-12){3}
//: {4}(34,31)(7,31)(7,10){5}
wire [31:0] w20;    //: /sn:0 {0}(-207,209)(-207,405){1}
//: {2}(-205,407)(-94,407)(-94,536)(194,536){3}
//: {4}(-209,407)(-218,407){5}
wire [31:0] w41;    //: /sn:0 {0}(-21,575)(194,575){1}
wire [31:0] w23;    //: /sn:0 /dp:17 {0}(-739,631)(-662,631)(-662,455)(-686,455){1}
//: {2}(-687,455)(-724,455){3}
//: {4}(-725,455)(-739,455){5}
//: {6}(-740,455)(-763,455){7}
//: {8}(-764,455)(-785,455){9}
//: {10}(-786,455)(-805,455){11}
//: {12}(-806,455)(-850,455){13}
//: {14}(-851,455)(-898,455){15}
//: {16}(-899,455)(-1232,455){17}
wire [4:0] w1;    //: /sn:0 {0}(-542,267)(-555,267){1}
//: {2}(-559,267)(-848,267){3}
//: {4}(-850,265)(-850,218){5}
//: {6}(-850,269)(-850,450){7}
//: {8}(-557,269)(-557,401)(-342,401){9}
wire [1:0] w25;    //: /sn:0 /dp:1 {0}(-52,314)(-52,-12){1}
wire [25:0] w35;    //: /sn:0 {0}(-739,498)(-739,490){1}
//: {2}(-737,488)(-653,488){3}
//: {4}(-739,486)(-739,459){5}
//: {6}(-741,488)(-1076,488)(-1076,432){7}
wire w8;    //: /sn:0 {0}(-1170,407)(-1170,402){1}
wire [31:0] w18;    //: /sn:0 {0}(-208,602)(-208,587){1}
//: {2}(-206,585)(-50,585){3}
//: {4}(-208,583)(-208,493){5}
//: {6}(-206,491)(-46,491)(-46,393)(64,393)(64,346)(686,346){7}
//: {8}(-208,489)(-208,439)(-218,439){9}
wire w30;    //: /sn:0 /dp:1 {0}(607,278)(595,278)(595,83)(-62,83){1}
//: {2}(-66,83)(-1473,83){3}
//: {4}(-1477,83)(-1524,83)(-1524,61){5}
//: {6}(-1475,85)(-1475,377)(-1424,377){7}
//: {8}(-64,85)(-64,284)(-254,284)(-254,365){9}
wire [15:0] w17;    //: /sn:0 {0}(-785,459)(-785,478)(-820,478)(-820,518){1}
//: {2}(-818,520)(-653,520){3}
//: {4}(-820,522)(-820,532)(-792,532){5}
//: {6}(-788,532)(-756,532){7}
//: {8}(-790,534)(-790,584)(-507,584)(-507,594){9}
wire [31:0] w22;    //: /sn:0 {0}(-1387,388)(-1387,461)(-1312,461)(-1312,458){1}
//: {2}(-1310,456)(-1302,456)(-1302,457)(-1290,457){3}
//: {4}(-1289,457)(-1267,457){5}
//: {6}(-1312,454)(-1312,362)(-1184,362){7}
wire [31:0] ReadData;    //: /sn:0 /dp:1 {0}(664,404)(700,404){1}
//: {2}(704,404)(712,404)(712,346)(702,346){3}
//: {4}(702,406)(702,426)(734,426){5}
wire [31:0] w53;    //: /sn:0 {0}(-1081,426)(-1081,399)(-1122,399)(-1122,255){1}
wire w57;    //: /sn:0 {0}(922,-12)(922,49){1}
//: {2}(920,51)(893,51)(893,15){3}
//: {4}(922,53)(922,483)(654,483)(654,467){5}
//: {6}(654,463)(654,431){7}
//: {8}(652,465)(616,465)(616,457){9}
wire [31:0] w2;    //: /sn:0 /dp:1 {0}(-1218,394)(-1184,394){1}
wire [2:0] w12;    //: /sn:0 {0}(7,360)(165,360)(165,392){1}
//: {2}(167,394)(258,394)(258,389){3}
//: {4}(165,396)(165,487)(222,487)(222,508){5}
wire [31:0] w10;    //: /sn:0 {0}(734,446)(702,446)(702,511)(522,511)(522,382)(503,382){1}
//: {2}(499,382)(382,382)(382,568)(256,568){3}
//: {4}(501,384)(501,417)(568,417)(568,409){5}
//: {6}(570,407)(601,407)(601,406)(629,406){7}
//: {8}(568,405)(568,363)(511,363)(511,326){9}
wire [4:0] w27;    //: /sn:0 {0}(-542,299)(-570,299){1}
//: {2}(-574,299)(-803,299){3}
//: {4}(-805,297)(-805,217){5}
//: {6}(-805,301)(-805,450){7}
//: {8}(-572,301)(-572,415)(-434,415){9}
//: {10}(-430,415)(-344,415){11}
//: {12}(-432,417)(-432,466)(-393,466){13}
wire [5:0] w13;    //: /sn:0 {0}(-617,-12)(-617,233){1}
//: {2}(-615,235)(-593,235){3}
//: {4}(-619,235)(-896,235){5}
//: {6}(-898,233)(-898,219){7}
//: {8}(-898,237)(-898,450){9}
wire [5:0] w52;    //: /sn:0 /dp:1 {0}(-1139,382)(-1139,442)(-1086,442)(-1086,432){1}
wire [31:0] w33;    //: /sn:0 /dp:1 {0}(856,581)(856,538)(778,538)(778,498){1}
//: {2}(778,494)(778,436)(763,436){3}
//: {4}(776,496)(-303,496)(-303,480){5}
wire [4:0] w5;    //: /sn:0 {0}(-542,331)(-578,331){1}
//: {2}(-582,331)(-761,331){3}
//: {4}(-763,329)(-763,218){5}
//: {6}(-763,333)(-763,450){7}
//: {8}(-580,333)(-580,446)(-393,446){9}
wire w29;    //: /sn:0 {0}(-439,-12)(-439,34){1}
//: {2}(-441,36)(-459,36)(-459,14){3}
//: {4}(-439,38)(-439,492)(-377,492)(-377,479){5}
wire [3:0] w9;    //: /sn:0 {0}(-662,434)(-662,439)(-643,439){1}
wire [31:0] w50;    //: /sn:0 {0}(-1089,316)(-1089,287)(-1102,287)(-1102,255){1}
wire [31:0] w39;    //: /sn:0 /dp:1 {0}(-1387,367)(-1387,192)(-1112,192)(-1112,226){1}
wire w26;    //: /sn:0 {0}(-485,-12)(-485,33){1}
//: {2}(-487,35)(-511,35)(-511,13){3}
//: {4}(-485,37)(-485,582)(-251,582)(-251,480){5}
//: enddecls

  //: switch g4 (w31) @(312,145) /sn:0 /R:3 /w:[ 5 ] /st:0
  led g8 (.I(w0));   //: @(-1270,565) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: joint g58 (w10) @(568, 407) /w:[ 6 8 -1 5 ]
  //: comment g37 /dolink:0 /link:"" @(-701,186) /sn:0 /R:3 /anc:1
  //: /line:"funct"
  //: /end
  led g13 (.I(w1));   //: @(-850,211) /sn:0 /anc:1 /w:[ 5 ] /type:1
  led g55 (.I(w26));   //: @(-511,6) /sn:0 /w:[ 3 ] /type:0
  bufif1 g139 (.Z(ReadData), .I(w18), .E(w45));   //: @(692,346) /sn:0 /w:[ 3 7 3 ]
  mux g76 (.I0(w27), .I1(w5), .S(w29), .Z(w46));   //: @(-377,456) /sn:0 /R:1 /w:[ 13 9 5 1 ] /ss:0 /do:0
  rom mRom (.A(w22), .D(w23), .OE(w4));   //: @(-1249,456) /sn:0 /w:[ 5 17 1 ]
  add g1 (.A(w2), .B(w22), .S(w7), .CI(w3), .CO(w8));   //: @(-1168,378) /sn:0 /R:1 /w:[ 1 7 0 1 1 ]
  register PC (.Q(w22), .D(w39), .EN(w11), .CLR(!w31), .CK(w30));   //: @(-1387,377) /sn:0 /w:[ 0 0 1 3 7 ]
  led g64 (.I(w21));   //: @(547,7) /sn:0 /w:[ 5 ] /type:0
  tran g11(.Z(w0), .I(w22[29:0]));   //: @(-1289,455) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  led g130 (.I(w12));   //: @(258,382) /sn:0 /w:[ 3 ] /type:3
  //: joint g121 (w28) @(36, 31) /w:[ -1 2 4 1 ]
  ALU g50 (.ALUop(w12), .B(w41), .A(w20), .Z(w19), .R(w10));   //: @(195, 509) /sz:(60, 101) /sn:0 /p:[ Ti0>5 Li0>1 Li1>3 Bo0<1 Ro0<3 ]
  led g28 (.I(w17));   //: @(-749,532) /sn:0 /R:3 /w:[ 7 ] /type:1
  //: joint g132 (w45) @(642, 330) /w:[ 2 1 -1 4 ]
  concat g113 (.I0(w35), .I1(w52), .Z(w53));   //: @(-1081,427) /sn:0 /R:1 /w:[ 7 1 0 ] /dr:0
  tran g19(.Z(w27), .I(w23[20:16]));   //: @(-805,453) /sn:0 /R:1 /w:[ 7 12 11 ] /ss:0
  //: comment g38 /dolink:0 /link:"" @(-735,541) /sn:0 /R:3
  //: /line:"address"
  //: /end
  //: dip g6 (w2) @(-1256,394) /sn:0 /R:1 /w:[ 0 ] /st:1
  CONTROL g53 (.op(w13), .Jump(w6), .Branch(w32), .RegDst(w29), .ALUsrc(w28), .RegWrite(w26), .ALUop(w25), .MemRead(w57), .MemWrite(w21), .MemToReg(w38));   //: @(-1662, -55) /sz:(2798, 42) /sn:0 /p:[ Bi0>0 Bo0<3 Bo1<5 Bo2<0 Bo3<3 Bo4<0 Bo5<1 Bo6<0 Bo7<3 Bo8<3 ]
  //: comment g75 /dolink:0 /link:"" @(-396,498) /sn:0
  //: /line:"RegDst"
  //: /line:"Seleciona "
  //: /line:"Reg Esc."
  //: /line:"rd -> R (1)"
  //: /line:"rt -> I (0)"
  //: /end
  //: supply0 g7 (w3) @(-1170,327) /sn:0 /R:2 /w:[ 0 ]
  //: joint g135 (w57) @(654, 465) /w:[ -1 6 8 5 ]
  //: comment g31 /dolink:0 /link:"" @(-1218,526) /sn:0 /R:3
  //: /line:"index"
  //: /end
  led g20 (.I(w5));   //: @(-763,211) /sn:0 /anc:1 /w:[ 5 ] /type:1
  //: joint g124 (w26) @(-485, 35) /w:[ -1 1 2 4 ]
  led g68 (.I(w33));   //: @(856,588) /sn:0 /R:2 /w:[ 0 ] /type:3
  Reg_32bits g39 (.Clock(w30), .Clear(w31), .R1(w1), .R2(w27), .Wr(w46), .Wd(w33), .RegWrite(w26), .D2(w18), .D1(w20));   //: @(-343, 366) /sz:(124, 113) /sn:0 /p:[ Ti0>9 Ti1>0 Li0>9 Li1>11 Li2>0 Bi0>5 Bi1>5 Ro0<9 Ro1<5 ]
  led g48 (.I(w18));   //: @(-208,609) /sn:0 /R:2 /w:[ 0 ] /type:3
  tran g29(.Z(w17), .I(w23[15:0]));   //: @(-785,453) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  tran g25(.Z(w15), .I(w23[5:0]));   //: @(-686,453) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:0
  tran g17(.Z(w13), .I(w23[31:26]));   //: @(-898,453) /sn:0 /R:1 /w:[ 9 16 15 ] /ss:0
  //: joint g52 (w18) @(-208, 585) /w:[ 2 4 -1 1 ]
  led g106 (.I(w35));   //: @(-646,488) /sn:0 /R:3 /w:[ 3 ] /type:3
  led g107 (.I(w17));   //: @(-646,520) /sn:0 /R:3 /w:[ 3 ] /type:3
  //: comment g83 /dolink:0 /link:"" @(244,212) /sn:0
  //: /line:"Branch"
  //: /line:"target"
  //: /end
  //: joint g100 (w13) @(-898, 235) /anc:1 /w:[ 5 6 -1 8 ]
  ram mRam (.A(w10), .D(ReadData), .WE(!w45), .OE(!w57), .CS(w36));   //: @(647,405) /sn:0 /delay:" 1 1 1 1 1 1 1" /w:[ 7 0 9 7 1 ]
  led g14 (.I(w13));   //: @(-898,212) /sn:0 /anc:1 /w:[ 7 ] /type:1
  led g47 (.I(w20));   //: @(-207,202) /sn:0 /w:[ 0 ] /type:3
  led g94 (.I(w13));   //: @(-586,235) /sn:0 /R:3 /w:[ 3 ] /type:3
  led g44 (.I(w32));   //: @(-905,17) /sn:0 /w:[ 7 ] /type:0
  //: joint g80 (w57) @(922, 51) /w:[ -1 1 2 4 ]
  led g84 (.I(w43));   //: @(236,305) /sn:0 /R:2 /w:[ 5 ] /type:3
  led g21 (.I(w14));   //: @(-724,210) /sn:0 /anc:1 /w:[ 5 ] /type:1
  //: joint g105 (w15) @(-686, 426) /w:[ 2 6 -1 1 ]
  tran g23(.Z(w14), .I(w23[10:6]));   //: @(-724,453) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:0
  //: joint g41 (w27) @(-432, 415) /w:[ 10 -1 9 12 ]
  //: joint g40 (w45) @(647, 369) /w:[ 6 5 -1 8 ]
  led g54 (.I(w10));   //: @(511,319) /sn:0 /w:[ 9 ] /type:3
  //: joint g93 (w37) @(-317, 671) /w:[ 2 -1 1 8 ]
  //: joint g123 (w29) @(-439, 36) /w:[ -1 1 2 4 ]
  //: joint g46 (w33) @(778, 496) /w:[ -1 2 4 1 ]
  led g26 (.I(w35));   //: @(-739,505) /sn:0 /R:2 /w:[ 0 ] /type:1
  //: supply0 g0 (w11) @(-1340,415) /sn:0 /w:[ 0 ]
  //: joint g90 (w38) @(832, 40) /w:[ -1 2 1 4 ]
  BEQ g82 (.PC(w7), .Btarget(w37), .Sum(w43));   //: @(106, 210) /sz:(81, 100) /sn:0 /p:[ Li0>7 Li1>7 Ro0<0 ]
  led g136 (.I(w23));   //: @(-746,631) /sn:0 /R:1 /w:[ 0 ] /type:2
  //: comment g128 /dolink:0 /link:"" @(-477,294) /sn:0
  //: /line:"R2"
  //: /end
  //: comment g33 /dolink:0 /link:"" @(-856,186) /sn:0 /R:3 /anc:1
  //: /line:"rs"
  //: /end
  //: comment g91 /dolink:0 /link:"" @(-1016,345) /sn:0 /R:2
  //: /line:"Branch-I"
  //: /end
  //: frame g49 @(-409,230) /sn:0 /wi:286 /ht:338 /tx:"BANC DE REGISTRES"
  //: comment g137 /dolink:0 /link:"" @(627,517) /sn:0
  //: /line:"D "
  //: /line:"(Read (1) de Lectura"
  //: /line:"(Write(1) de Escritura"
  //: /end
  //: comment g61 /dolink:0 /link:"" @(770,361) /sn:0
  //: /line:"MemtoReg"
  //: /end
  //: joint g86 (w37) @(-76, 565) /w:[ 4 6 -1 3 ]
  mux g3 (.I0(w50), .I1(w53), .S(w6), .Z(w39));   //: @(-1112,239) /sn:0 /R:2 /w:[ 1 1 5 1 ] /ss:0 /do:0
  //: joint g51 (w20) @(-207, 407) /w:[ 2 1 4 -1 ]
  //: comment g34 /dolink:0 /link:"" @(-809,185) /sn:0 /R:3 /anc:1
  //: /line:"rt"
  //: /end
  mux g89 (.I0(w7), .I1(w43), .S(w34), .Z(w50));   //: @(-1089,329) /sn:0 /R:2 /w:[ 5 3 0 0 ] /ss:0 /do:0
  led g2 (.I(w45));   //: @(674,351) /sn:0 /w:[ 7 ] /type:0
  //: joint g65 (w13) @(-617, 235) /w:[ 2 1 4 -1 ]
  //: joint g77 (w5) @(-580, 331) /w:[ 1 -1 2 8 ]
  //: comment g110 /dolink:0 /link:"" @(-1022,248) /sn:0
  //: /line:"Branch-J"
  //: /end
  mux g59 (.I0(w10), .I1(ReadData), .S(w38), .Z(w33));   //: @(750,436) /sn:0 /R:1 /w:[ 0 5 5 3 ] /ss:0 /do:0
  //: joint g72 (w17) @(-790, 532) /w:[ 6 -1 5 8 ]
  led g98 (.I(w14));   //: @(-641,394) /sn:0 /R:3 /w:[ 3 ] /type:3
  led g99 (.I(w9));   //: @(-636,439) /sn:0 /R:3 /w:[ 1 ] /type:3
  led g96 (.I(w27));   //: @(-535,299) /sn:0 /R:3 /w:[ 0 ] /type:3
  led g16 (.I(w6));   //: @(-976,16) /sn:0 /w:[ 0 ] /type:0
  //: joint g122 (w1) @(-557, 267) /w:[ 1 -1 2 8 ]
  //: joint g103 (w5) @(-763, 331) /w:[ 3 4 -1 6 ]
  SignExtend16to32bits g78 (.Adr16(w17), .Adr32(w37));   //: @(-588, 595) /sz:(156, 60) /sn:0 /p:[ Ti0>9 Bo0<0 ]
  //: supply0 g10 (w4) @(-1149,529) /sn:0 /w:[ 0 ]
  //: joint g87 (w30) @(-1475, 83) /w:[ 3 -1 4 6 ]
  //: comment g129 /dolink:0 /link:"" @(-476,327) /sn:0
  //: /line:"Rd"
  //: /end
  //: comment g32 /dolink:0 /link:"" @(-825,-7) /sn:0 /R:3
  //: /line:"clear"
  //: /end
  tran g27(.Z(w35), .I(w23[25:0]));   //: @(-739,453) /sn:0 /R:1 /w:[ 5 6 5 ] /ss:1
  //: joint g102 (w27) @(-805, 299) /anc:1 /w:[ 3 4 -1 6 ]
  mux g69 (.I0(w18), .I1(w37), .S(w28), .Z(w41));   //: @(-34,575) /sn:0 /R:1 /w:[ 3 5 0 0 ] /ss:0 /do:0
  //: comment g57 /dolink:0 /link:"" @(196,418) /sn:0
  //: /line:"0000 (0) -> AND (A&b)"
  //: /line:"0001 (1) -> OR 	 (AoB)"
  //: /line:"0010 (2) -> ADD	 (A+B)"
  //: /line:"0110 (6) -> SUB (A-B)"
  //: /line:"0111 (7) -> SLT	 (A<B)"
  //: /end
  clock g9 (.Z(w30));   //: @(-1521,49) /sn:0 /R:3 /anc:1 /w:[ 5 ] /omega:566 /phi:0 /duty:50
  //: joint g119 (w21) @(570, 35) /w:[ -1 2 4 1 ]
  //: comment g71 /dolink:0 /link:"" @(-31,612) /sn:0
  //: /line:"ALUsrc"
  //: /line:"Selecion: "
  //: /line:"Operand 2 "
  //: /line:"BancoReg	(0)"
  //: /line:"Instrucc	(1)"
  //: /end
  led g15 (.I(w27));   //: @(-805,210) /sn:0 /anc:1 /w:[ 5 ] /type:1
  //: joint g131 (w12) @(165, 394) /w:[ 2 1 -1 4 ]
  //: comment g127 /dolink:0 /link:"" @(-478,261) /sn:0
  //: /line:"R1"
  //: /end
  tran g67(.Z(w9), .I(w15[3:0]));   //: @(-662,424) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  and g43 (.I0(w19), .I1(w32), .Z(w34));   //: @(-993,375) /sn:0 /R:2 /w:[ 0 0 1 ]
  //: joint g88 (w7) @(-1097, 378) /w:[ 4 6 3 -1 ]
  //: comment g73 /dolink:0 /link:"" @(-1395,370) /sn:0
  //: /line:"PC"
  //: /end
  //: joint g104 (w14) @(-724, 394) /w:[ 2 4 -1 1 ]
  led g62 (.I(w29));   //: @(-459,7) /sn:0 /w:[ 3 ] /type:0
  //: supply0 g138 (w36) @(635,476) /sn:0 /w:[ 0 ]
  //: joint g42 (w30) @(-64, 83) /w:[ 1 -1 2 8 ]
  led g63 (.I(w28));   //: @(7,3) /sn:0 /w:[ 5 ] /type:0
  //: joint g109 (w35) @(-739, 488) /w:[ 2 4 6 1 ]
  led g74 (.I(w57));   //: @(893,8) /sn:0 /w:[ 3 ] /type:0
  //: joint g5 (w22) @(-1312, 456) /w:[ 2 6 -1 1 ]
  //: joint g56 (ReadData) @(702, 404) /w:[ 2 -1 1 4 ]
  //: joint g133 (w10) @(501, 382) /w:[ 1 -1 2 4 ]
  and g79 (.I0(w30), .I1(w21), .Z(w45));   //: @(618,281) /sn:0 /w:[ 0 0 0 ]
  led g95 (.I(w1));   //: @(-535,267) /sn:0 /R:3 /w:[ 0 ] /type:3
  ALUctr g117 (.SelOp(w25), .funct(w15), .Oop(w12));   //: @(-109, 315) /sz:(115, 64) /sn:0 /p:[ Ti0>0 Li0>5 Ro0<0 ]
  //: comment g36 /dolink:0 /link:"" @(-741,185) /sn:0 /R:3 /anc:1
  //: /line:"shamt"
  //: /end
  led g24 (.I(w15));   //: @(-686,210) /sn:0 /anc:1 /w:[ 7 ] /type:1
  //: joint g85 (w43) @(236, 227) /w:[ -1 2 1 4 ]
  led g92 (.I(w37));   //: @(-317,697) /sn:0 /R:2 /w:[ 9 ] /type:3
  //: comment g144 /dolink:0 /link:"" @(682,308) /sn:0
  //: /line:"Leer o Escribir"
  //: /end
  //: joint g125 (w32) @(-926, 45) /w:[ 2 4 6 1 ]
  //: joint g101 (w1) @(-850, 267) /anc:1 /w:[ 3 4 -1 6 ]
  //: joint g60 (w18) @(-208, 491) /w:[ 6 8 -1 5 ]
  //: frame g81 @(70,98) /sn:0 /wi:299 /ht:249 /tx:"ALU-I"
  led g70 (.I(w38));   //: @(790,10) /sn:0 /w:[ 0 ] /type:0
  //: frame g45 @(71,404) /sn:0 /wi:298 /ht:344 /tx:"ALU-R"
  //: joint g126 (w6) @(-1003, 43) /w:[ 1 2 -1 4 ]
  //: comment g35 /dolink:0 /link:"" @(-768,186) /sn:0 /R:3 /anc:1
  //: /line:"rd"
  //: /end
  tran g22(.Z(w5), .I(w23[15:11]));   //: @(-763,453) /sn:0 /R:1 /w:[ 7 8 7 ] /ss:0
  //: joint g120 (w27) @(-572, 299) /w:[ 1 -1 2 8 ]
  tran g114(.Z(w52), .I(w7[31:26]));   //: @(-1139,376) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: frame g66 @(400,222) /sn:0 /wi:479 /ht:341 /tx:"DATA MEMORY"
  led g97 (.I(w5));   //: @(-535,331) /sn:0 /R:3 /w:[ 0 ] /type:3
  tran g18(.Z(w1), .I(w23[25:21]));   //: @(-850,453) /sn:0 /R:1 /w:[ 7 14 13 ] /ss:0
  //: frame g12 @(-1463,174) /sn:0 /wi:517 /ht:427 /tx:"FETCH"
  //: comment g30 /dolink:0 /link:"" @(-901,185) /sn:0 /R:3 /anc:1
  //: /line:"op"
  //: /end
  //: joint g108 (w17) @(-820, 520) /w:[ 2 1 -1 4 ]
  //: joint g118 (w31) @(-808, 60) /w:[ 1 -1 2 4 ]
  led g134 (.I(w57));   //: @(616,450) /sn:0 /w:[ 9 ] /type:0

endmodule

module Intruction_Memory(Instruction, Read_Address);
//: interface  /sz:(40, 40) /bd:[ Li0>Read_Address[7:0](10/40) Li1>Read_Address[7:0](10/40) Ro0<Instruction[7:0](24/40) Ro1<Instruction[7:0](24/40) ]
input Read_Address;    //: /sn:0 {0}(148,118)(158,118){1}
output Instruction;    //: /sn:0 /dp:1 {0}(467,116)(477,116){1}
//: enddecls

  //: output g1 (Instruction) @(474,116) /sn:0 /w:[ 1 ]
  //: input g0 (Read_Address) @(146,118) /sn:0 /w:[ 0 ]

endmodule

module ALUctr(Oop, SelOp, funct);
//: interface  /sz:(40, 40) /bd:[ ]
input [1:0] SelOp;    //: /sn:0 /dp:1 {0}(215,204)(215,233){1}
//: {2}(215,234)(215,267){3}
//: {4}(215,268)(215,276){5}
input [5:0] funct;    //: /sn:0 {0}(175,249)(175,281){1}
//: {2}(175,282)(175,315){3}
//: {4}(175,316)(175,355){5}
//: {6}(175,356)(175,369){7}
//: {8}(175,370)(175,380){9}
output [2:0] Oop;    //: /sn:0 /dp:1 {0}(535,319)(608,319){1}
wire w7;    //: /sn:0 /dp:1 {0}(343,286)(198,286)(198,356)(179,356){1}
wire w16;    //: /sn:0 /dp:1 {0}(351,370)(179,370){1}
wire w14;    //: /sn:0 {0}(421,282)(452,282)(452,309)(529,309){1}
wire w4;    //: /sn:0 /dp:1 {0}(529,329)(452,329)(452,349)(442,349){1}
wire w18;    //: /sn:0 {0}(219,234)(365,234)(365,268)(381,268)(381,279)(400,279){1}
wire w8;    //: /sn:0 {0}(424,319)(529,319){1}
wire w2;    //: /sn:0 {0}(372,368)(394,368)(394,351)(421,351){1}
wire w11;    //: /sn:0 {0}(364,284)(400,284){1}
wire w12;    //: /sn:0 {0}(219,268)(313,268)(313,280){1}
//: {2}(315,282)(325,282)(325,281)(343,281){3}
//: {4}(313,284)(313,335)(391,335){5}
//: {6}(393,333)(393,321)(403,321){7}
//: {8}(393,337)(393,346)(421,346){9}
wire w10;    //: /sn:0 /dp:1 {0}(403,316)(179,316){1}
wire w9;    //: /sn:0 {0}(179,282)(273,282)(273,365)(351,365){1}
//: enddecls

  and g4 (.I0(w12), .I1(w2), .Z(w4));   //: @(432,349) /sn:0 /w:[ 9 1 1 ]
  tran g8(.Z(w16), .I(funct[0]));   //: @(173,370) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  //: joint g13 (w12) @(313, 282) /w:[ 2 1 -1 4 ]
  or g3 (.I0(w9), .I1(w16), .Z(w2));   //: @(362,368) /sn:0 /w:[ 1 0 0 ]
  //: output g2 (Oop) @(605,319) /sn:0 /w:[ 1 ]
  //: input g1 (SelOp) @(215,202) /sn:0 /R:3 /w:[ 0 ]
  tran g11(.Z(w10), .I(funct[2]));   //: @(173,316) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  tran g16(.Z(w9), .I(funct[3]));   //: @(173,282) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  concat g10 (.I0(w4), .I1(w8), .I2(w14), .Z(Oop));   //: @(534,319) /sn:0 /w:[ 0 1 1 0 ] /dr:0
  and g6 (.I0(w12), .I1(w7), .Z(w11));   //: @(354,284) /sn:0 /w:[ 3 0 0 ]
  or g7 (.I0(w18), .I1(w11), .Z(w14));   //: @(411,282) /sn:0 /w:[ 1 1 0 ]
  tran g9(.Z(w7), .I(funct[1]));   //: @(173,356) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  tran g15(.Z(w12), .I(SelOp[1]));   //: @(213,268) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  or g5 (.I0(!w10), .I1(!w12), .Z(w8));   //: @(414,319) /sn:0 /w:[ 0 7 0 ]
  tran g14(.Z(w18), .I(SelOp[0]));   //: @(213,234) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g0 (funct) @(175,247) /sn:0 /R:3 /w:[ 0 ]
  //: joint g12 (w12) @(393, 335) /w:[ -1 6 5 8 ]

endmodule
