//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(477,287)(273,287)(273,216){1}
wire w7;    //: /sn:0 {0}(292,192)(334,192){1}
wire w16;    //: /sn:0 {0}(445,128)(445,174){1}
wire [7:0] w4;    //: /sn:0 {0}(72,110)(72,124)(193,124){1}
//: {2}(194,124)(276,124){3}
//: {4}(277,124)(360,124){5}
//: {6}(361,124)(444,124){7}
//: {8}(445,124)(583,124){9}
wire w15;    //: /sn:0 {0}(361,128)(361,174){1}
wire w3;    //: /sn:0 {0}(194,128)(194,174){1}
wire w0;    //: /sn:0 {0}(183,68)(183,174){1}
wire [4:0] w21;    //: /sn:0 /dp:1 {0}(483,287)(576,287){1}
wire [3:0] w24;    //: /sn:0 /dp:9 {0}(576,64)(434,64){1}
//: {2}(433,64)(350,64){3}
//: {4}(349,64)(266,64){5}
//: {6}(265,64)(183,64){7}
//: {8}(182,64)(72,64)(72,59){9}
wire w20;    //: /sn:0 /dp:1 {0}(477,297)(357,297)(357,216){1}
wire w1;    //: /sn:0 {0}(266,68)(266,174){1}
wire w18;    //: /sn:0 /dp:1 {0}(477,307)(441,307)(441,216){1}
wire w8;    //: /sn:0 {0}(209,192)(250,192){1}
wire w22;    //: /sn:0 {0}(477,277)(190,277)(190,216){1}
wire w11;    //: /sn:0 {0}(277,128)(277,174){1}
wire w12;    //: /sn:0 {0}(434,68)(434,174){1}
wire w10;    //: /sn:0 /dp:1 {0}(477,267)(120,267)(120,194){1}
//: {2}(122,192)(167,192){3}
//: {4}(118,192)(91,192)(91,180){5}
wire w13;    //: /sn:0 {0}(376,192)(418,192){1}
wire w5;    //: /sn:0 {0}(499,192)(460,192){1}
wire w9;    //: /sn:0 {0}(350,68)(350,174){1}
//: enddecls

  led g8 (.I(w10));   //: @(91,173) /sn:0 /w:[ 5 ] /type:0
  SFA g4 (.B(w11), .A(w1), .Ci(w7), .Co(w8), .S(w6));   //: @(251, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  tran g13(.Z(w9), .I(w24[1]));   //: @(350,62) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g3(.Z(w0), .I(w24[3]));   //: @(183,62) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  led g2 (.I(w21));   //: @(583,287) /sn:0 /R:3 /w:[ 1 ] /type:3
  //: dip g1 (w24) @(72,49) /sn:0 /w:[ 9 ] /st:9
  tran g16(.Z(w16), .I(w4[0]));   //: @(445,122) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g11(.Z(w1), .I(w24[2]));   //: @(266,62) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g10(.Z(w3), .I(w4[3]));   //: @(194,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g19 (w10) @(120, 192) /w:[ 2 -1 4 1 ]
  SFA g6 (.B(w16), .A(w12), .Ci(w5), .Co(w13), .S(w18));   //: @(419, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: dip g9 (w4) @(72,100) /sn:0 /w:[ 0 ] /st:0
  concat g7 (.I0(w18), .I1(w20), .I2(w6), .I3(w22), .I4(w10), .Z(w21));   //: @(482,287) /sn:0 /w:[ 0 0 0 0 0 0 ] /dr:0
  tran g15(.Z(w15), .I(w4[1]));   //: @(361,122) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: switch g17 (w5) @(517,192) /sn:0 /R:2 /w:[ 0 ] /st:1
  tran g14(.Z(w12), .I(w24[0]));   //: @(434,62) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  SFA g5 (.B(w15), .A(w9), .Ci(w13), .Co(w7), .S(w20));   //: @(335, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  SFA g0 (.B(w3), .A(w0), .Ci(w8), .Co(w10), .S(w22));   //: @(168, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<3 Bo0<1 ]
  tran g12(.Z(w11), .I(w4[2]));   //: @(277,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module SFA(S, Ci, B, A, Co);
//: interface  /sz:(40, 40) /bd:[ Ti0>A(15/40) Ti1>B(26/40) Ri0>Ci(17/40) Lo0<Co(17/40) Bo0<S(22/40) ]
input B;    //: /sn:0 {0}(66,121)(105,121){1}
//: {2}(109,121)(149,121)(149,103)(157,103){3}
//: {4}(107,123)(107,193)(163,193){5}
input A;    //: /sn:0 /dp:1 {0}(157,98)(99,98)(99,102){1}
//: {2}(97,104)(65,104){3}
//: {4}(99,106)(99,188)(163,188){5}
output Co;    //: /sn:0 {0}(288,178)(249,178){1}
input Ci;    //: /sn:0 {0}(67,141)(132,141){1}
//: {2}(136,141)(212,141)(212,127)(220,127){3}
//: {4}(134,143)(134,162)(164,162){5}
output S;    //: /sn:0 {0}(286,125)(241,125){1}
wire w8;    //: /sn:0 {0}(184,191)(218,191)(218,180)(228,180){1}
wire w2;    //: /sn:0 {0}(178,101)(190,101){1}
//: {2}(194,101)(210,101)(210,122)(220,122){3}
//: {4}(192,103)(192,132)(155,132)(155,167)(164,167){5}
wire w5;    //: /sn:0 {0}(185,165)(218,165)(218,175)(228,175){1}
//: enddecls

  //: joint g8 (A) @(99, 104) /w:[ -1 1 2 4 ]
  and g4 (.I0(Ci), .I1(w2), .Z(w5));   //: @(175,165) /sn:0 /w:[ 5 5 0 ]
  //: output g13 (S) @(283,125) /sn:0 /w:[ 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(168,101) /sn:0 /w:[ 0 3 0 ]
  //: input g2 (Ci) @(65,141) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(64,121) /sn:0 /w:[ 0 ]
  //: joint g11 (w2) @(192, 101) /w:[ 2 -1 1 4 ]
  //: joint g10 (Ci) @(134, 141) /w:[ 2 -1 1 4 ]
  or g6 (.I0(w5), .I1(w8), .Z(Co));   //: @(239,178) /sn:0 /w:[ 1 1 1 ]
  //: joint g9 (B) @(107, 121) /w:[ 2 -1 1 4 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(231,125) /sn:0 /w:[ 3 3 1 ]
  and g5 (.I0(A), .I1(B), .Z(w8));   //: @(174,191) /sn:0 /w:[ 5 5 0 ]
  //: input g0 (A) @(63,104) /sn:0 /w:[ 3 ]
  //: output g12 (Co) @(285,178) /sn:0 /w:[ 0 ]

endmodule
