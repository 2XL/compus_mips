//: version "1.8.7"

module CaLoA(cf, p, g, ci);
//: interface  /sz:(40, 40) /bd:[ Ti0>g(28/40) Ti1>p(10/40) Ri0>ci(22/40) Lo0<cf(20/40) ]
input p;    //: /sn:0 {0}(105,123)(163,123)(163,134)(173,134){1}
output cf;    //: /sn:0 /dp:1 {0}(261,99)(319,99){1}
input ci;    //: /sn:0 {0}(109,150)(163,150)(163,139)(173,139){1}
input g;    //: /sn:0 {0}(107,87)(230,87)(230,96)(240,96){1}
wire w2;    //: /sn:0 {0}(194,137)(230,137)(230,101)(240,101){1}
//: enddecls

  xor g4 (.I0(p), .I1(ci), .Z(w2));   //: @(184,137) /sn:0 /w:[ 1 1 0 ]
  //: output g3 (cf) @(316,99) /sn:0 /w:[ 1 ]
  //: input g2 (p) @(103,123) /sn:0 /w:[ 0 ]
  //: input g1 (g) @(105,87) /sn:0 /w:[ 0 ]
  and g5 (.I0(g), .I1(w2), .Z(cf));   //: @(251,99) /sn:0 /w:[ 1 1 0 ]
  //: input g0 (ci) @(107,150) /sn:0 /w:[ 0 ]

endmodule

module Carrylookahead_logic(p3, c3, g3, c2, c1, p1, g0, c4, g2, g1, p2, c0, p0);
//: interface  /sz:(379, 40) /bd:[ Ti0>g0(321/379) Ti1>p0(311/379) Ti2>g1(233/379) Ti3>p1(225/379) Ti4>g2(144/379) Ti5>p2(135/379) Ti6>g3(58/379) Ti7>p3(50/379) Ri0>c0(24/40) To0<c3(95/379) To1<c2(182/379) To2<c1(272/379) Lo0<c4(20/40) ]
input g3;    //: /sn:0 {0}(179,35)(179,120){1}
input g2;    //: /sn:0 {0}(243,35)(243,82)(242,82)(242,122){1}
input c0;    //: /sn:0 {0}(64,-33)(509,-33)(509,149)(441,149){1}
input g1;    //: /sn:0 {0}(327,35)(327,88)(329,88)(329,124){1}
output c4;    //: /sn:0 {0}(150,141)(30,141){1}
output c1;    //: /sn:0 {0}(38,-16)(379,-16)(379,145){1}
//: {2}(381,147)(399,147){3}
//: {4}(377,147)(360,147){5}
input p3;    //: /sn:0 {0}(158,35)(158,82)(161,82)(161,120){1}
input p2;    //: /sn:0 {0}(260,35)(260,122){1}
output c3;    //: /sn:0 {0}(38,15)(209,15)(209,141){1}
//: {2}(211,143)(231,143){3}
//: {4}(207,143)(192,143){5}
input p1;    //: /sn:0 {0}(343,34)(343,87)(347,87)(347,124){1}
output c2;    //: /sn:0 {0}(69,0)(298,0)(298,143){1}
//: {2}(300,145)(318,145){3}
//: {4}(296,145)(273,145){5}
input p0;    //: /sn:0 {0}(412,41)(412,90)(410,90)(410,126){1}
input g0;    //: /sn:0 {0}(429,40)(429,94)(428,94)(428,126){1}
//: enddecls

  CaLoA g4 (.g(g3), .p(p3), .ci(c3), .cf(c4));   //: @(151, 121) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<0 ]
  //: input g8 (p3) @(158,33) /sn:0 /R:3 /w:[ 0 ]
  //: output g3 (c3) @(41,15) /sn:0 /R:2 /w:[ 0 ]
  //: input g13 (g3) @(179,33) /sn:0 /R:3 /w:[ 0 ]
  //: output g2 (c2) @(72,0) /sn:0 /R:2 /w:[ 0 ]
  //: output g1 (c1) @(41,-16) /sn:0 /R:2 /w:[ 0 ]
  //: joint g11 (c2) @(298, 145) /w:[ 2 1 4 -1 ]
  //: input g16 (p1) @(343,32) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (c1) @(379, 147) /w:[ 2 1 4 -1 ]
  //: input g19 (g0) @(429,38) /sn:0 /R:3 /w:[ 0 ]
  CaLoA g6 (.g(p1), .p(g1), .ci(c1), .cf(c2));   //: @(319, 125) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<3 ]
  CaLoA g7 (.g(g0), .p(p0), .ci(c0), .cf(c1));   //: @(400, 127) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<3 ]
  //: output g9 (c4) @(33,141) /sn:0 /R:2 /w:[ 1 ]
  //: input g15 (g2) @(243,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g17 (g1) @(327,33) /sn:0 /R:3 /w:[ 0 ]
  CaLoA g5 (.g(p2), .p(g2), .ci(c2), .cf(c3));   //: @(232, 123) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>5 Lo0<3 ]
  //: input g14 (p2) @(260,33) /sn:0 /R:3 /w:[ 0 ]
  //: input g0 (c0) @(62,-33) /sn:0 /w:[ 0 ]
  //: joint g12 (c3) @(209, 143) /w:[ 2 1 4 -1 ]
  //: input g18 (p0) @(412,39) /sn:0 /R:3 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(266,20)(266,155){1}
wire w7;    //: /sn:0 {0}(279,68)(279,155){1}
wire w19;    //: /sn:0 {0}(456,68)(456,156){1}
wire w4;    //: /sn:0 /dp:1 {0}(197,197)(197,376)(487,376){1}
wire w38;    //: /sn:0 {0}(353,197)(353,275)(357,275)(357,285){1}
wire w0;    //: /sn:0 {0}(180,20)(180,155){1}
wire w3;    //: /sn:0 {0}(314,285)(314,220)(308,220)(308,175)(293,175){1}
wire [3:0] w24;    //: /sn:0 {0}(82,16)(179,16){1}
//: {2}(180,16)(265,16){3}
//: {4}(266,16)(354,16){5}
//: {6}(355,16)(442,16){7}
//: {8}(443,16)(517,16){9}
wire w23;    //: /sn:0 {0}(460,198)(460,406)(487,406){1}
wire w20;    //: /sn:0 {0}(487,366)(93,366)(93,254)(115,254){1}
//: {2}(117,252)(117,217){3}
//: {4}(117,256)(117,306)(131,306){5}
wire w36;    //: /sn:0 {0}(274,197)(274,275)(276,275)(276,285){1}
wire w41;    //: /sn:0 {0}(441,198)(441,275)(443,275)(443,285){1}
wire w1;    //: /sn:0 {0}(193,68)(193,155){1}
wire [3:0] w25;    //: /sn:0 {0}(80,64)(192,64){1}
//: {2}(193,64)(278,64){3}
//: {4}(279,64)(367,64){5}
//: {6}(368,64)(455,64){7}
//: {8}(456,64)(517,64){9}
wire w18;    //: /sn:0 {0}(443,20)(443,156){1}
wire w35;    //: /sn:0 {0}(264,197)(264,275)(267,275)(267,285){1}
wire w8;    //: /sn:0 {0}(190,285)(190,226)(188,226)(188,197){1}
wire w17;    //: /sn:0 {0}(372,197)(372,396)(487,396){1}
wire w12;    //: /sn:0 {0}(355,20)(355,155){1}
wire w11;    //: /sn:0 /dp:1 {0}(283,197)(283,386)(487,386){1}
wire w2;    //: /sn:0 {0}(227,285)(227,175)(207,175){1}
wire w13;    //: /sn:0 {0}(368,68)(368,155){1}
wire [4:0] w33;    //: /sn:0 /dp:1 {0}(493,386)(555,386)(555,363){1}
wire w5;    //: /sn:0 {0}(404,285)(404,223)(398,223)(398,175)(382,175){1}
wire w42;    //: /sn:0 {0}(451,198)(451,275)(453,275)(453,285){1}
wire w9;    //: /sn:0 {0}(182,285)(182,225)(178,225)(178,197){1}
wire w26;    //: /sn:0 {0}(561,176)(533,176){1}
//: {2}(529,176)(470,176){3}
//: {4}(531,178)(531,310)(512,310){5}
wire w39;    //: /sn:0 {0}(363,197)(363,275)(365,275)(365,285){1}
//: enddecls

  tran g8(.Z(w12), .I(w24[1]));   //: @(355,14) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: dip g4 (w24) @(44,16) /sn:0 /R:1 /w:[ 0 ] /st:0
  tran g13(.Z(w1), .I(w25[3]));   //: @(193,62) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  S_CLA g3 (.B(w19), .A(w18), .C(w26), .S(w23), .G(w42), .P(w41));   //: @(429, 157) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<0 Bo1<0 Bo2<0 ]
  S_CLA g2 (.B(w13), .A(w12), .C(w5), .S(w17), .G(w39), .P(w38));   //: @(341, 156) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  S_CLA g1 (.B(w7), .A(w6), .C(w3), .S(w11), .G(w36), .P(w35));   //: @(252, 156) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  Carrylookahead_logic g16 (.p3(w9), .g3(w8), .p2(w35), .g2(w36), .p1(w38), .g1(w39), .p0(w41), .g0(w42), .c0(w26), .c1(w5), .c2(w3), .c3(w2), .c4(w20));   //: @(132, 286) /sz:(379, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<0 To1<0 To2<0 Lo0<5 ]
  tran g11(.Z(w19), .I(w25[0]));   //: @(456,62) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g10(.Z(w13), .I(w25[1]));   //: @(368,62) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  led g28 (.I(w20));   //: @(117,210) /sn:0 /w:[ 3 ] /type:0
  led g32 (.I(w33));   //: @(555,356) /sn:0 /w:[ 1 ] /type:3
  tran g6(.Z(w0), .I(w24[3]));   //: @(180,14) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g9(.Z(w18), .I(w24[0]));   //: @(443,14) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g7(.Z(w6), .I(w24[2]));   //: @(266,14) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g15 (w26) @(531, 176) /w:[ 1 -1 2 4 ]
  //: joint g17 (w20) @(117, 254) /w:[ -1 2 1 4 ]
  //: switch g14 (w26) @(579,176) /sn:0 /R:2 /w:[ 0 ] /st:0
  //: dip g5 (w25) @(42,64) /sn:0 /R:1 /w:[ 0 ] /st:0
  S_CLA g0 (.B(w1), .A(w0), .C(w2), .S(w4), .G(w8), .P(w9));   //: @(166, 156) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  tran g12(.Z(w7), .I(w25[2]));   //: @(279,62) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  concat g30 (.I0(w23), .I1(w17), .I2(w11), .I3(w4), .I4(w20), .Z(w33));   //: @(492,386) /sn:0 /w:[ 1 1 1 1 0 0 ] /dr:0

endmodule

module S_CLA(A, P, C, S, G, B);
//: interface  /sz:(40, 40) /bd:[ Ti0>A(14/40) Ti1>B(27/40) Ri0>C(19/40) Bo0<P(12/40) Bo1<G(22/40) Bo2<S(31/40) ]
input B;    //: /sn:0 {0}(-293,-95)(-250,-95){1}
//: {2}(-246,-95)(-223,-95)(-223,-105)(-149,-105){3}
//: {4}(-248,-93)(-248,-74){5}
//: {6}(-246,-72)(-35,-72){7}
//: {8}(-248,-70)(-248,-34)(-36,-34){9}
input A;    //: /sn:0 /dp:1 {0}(-149,-110)(-222,-110)(-222,-119)(-269,-119){1}
//: {2}(-273,-119)(-294,-119){3}
//: {4}(-271,-117)(-271,-69){5}
//: {6}(-269,-67)(-35,-67){7}
//: {8}(-271,-65)(-271,-29)(-36,-29){9}
output G;    //: /sn:0 /dp:1 {0}(-15,-31)(73,-31){1}
output P;    //: /sn:0 {0}(73,-69)(-14,-69){1}
input C;    //: /sn:0 {0}(-293,-80)(-62,-80)(-62,-120)(-37,-120){1}
output S;    //: /sn:0 /dp:1 {0}(-16,-122)(73,-122){1}
wire w3;    //: /sn:0 /dp:1 {0}(-37,-125)(-76,-125)(-76,-107)(-128,-107){1}
//: enddecls

  //: input g4 (A) @(-296,-119) /sn:0 /w:[ 3 ]
  //: output g8 (P) @(70,-69) /sn:0 /w:[ 0 ]
  and g3 (.I0(B), .I1(A), .Z(G));   //: @(-25,-31) /sn:0 /w:[ 9 9 0 ]
  //: joint g13 (B) @(-248, -72) /w:[ 6 5 -1 8 ]
  or g2 (.I0(B), .I1(A), .Z(P));   //: @(-24,-69) /sn:0 /w:[ 7 7 1 ]
  xor g1 (.I0(w3), .I1(C), .Z(S));   //: @(-26,-122) /sn:0 /w:[ 0 1 0 ]
  //: joint g11 (A) @(-271, -67) /w:[ 6 5 -1 8 ]
  //: joint g10 (A) @(-271, -119) /w:[ 1 -1 2 4 ]
  //: input g6 (C) @(-295,-80) /sn:0 /w:[ 0 ]
  //: output g7 (S) @(70,-122) /sn:0 /w:[ 1 ]
  //: output g9 (G) @(70,-31) /sn:0 /w:[ 1 ]
  //: input g5 (B) @(-295,-95) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(w3));   //: @(-138,-107) /sn:0 /w:[ 0 3 1 ]
  //: joint g12 (B) @(-248, -95) /w:[ 2 -1 1 4 ]

endmodule
