//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(-90,46)(-90,54)(-87,54)(-87,61){1}
wire w96;    //: /sn:0 /dp:1 {0}(-327,728)(-327,796)(429,796){1}
wire w7;    //: /sn:0 {0}(-85,82)(-85,175)(70,175)(70,242){1}
wire w99;    //: /sn:0 {0}(-485,708)(-349,708){1}
wire w61;    //: /sn:0 {0}(18,737)(18,816)(429,816){1}
wire w16;    //: /sn:0 {0}(-273,505)(-273,595)(-159,595)(-159,688){1}
wire w56;    //: /sn:0 {0}(-327,285)(-452,285)(-452,465){1}
wire w14;    //: /sn:0 {0}(-123,101)(-123,184){1}
wire [7:0] w19;    //: /sn:0 /dp:1 {0}(536,81)(536,811)(435,811){1}
wire w89;    //: /sn:0 /dp:1 {0}(-130,708)(-18,708)(-18,713)(-8,713){1}
wire w15;    //: /sn:0 {0}(-279,101)(-279,119)(-277,119)(-277,160){1}
wire w4;    //: /sn:0 {0}(-82,61)(-82,21){1}
//: {2}(-80,19)(128,19){3}
//: {4}(132,19)(285,19){5}
//: {6}(289,19)(379,19){7}
//: {8}(287,21)(287,31)(286,31)(286,64){9}
//: {10}(130,21)(130,60){11}
//: {12}(-84,19)(-160,19){13}
//: {14}(-164,19)(-596,19){15}
//: {16}(-162,21)(-162,59){17}
wire w38;    //: /sn:0 {0}(429,776)(-561,776)(-561,709)(-527,709){1}
wire w51;    //: /sn:0 {0}(-430,542)(-430,594)(-433,594)(-433,638){1}
wire w97;    //: /sn:0 /dp:1 {0}(-498,687)(-498,669)(-431,669)(-431,659){1}
wire w0;    //: /sn:0 {0}(381,130)(245,130){1}
//: {2}(241,130)(88,130){3}
//: {4}(84,130)(-116,130){5}
//: {6}(-120,130)(-270,130){7}
//: {8}(-274,130)(-596,130){9}
//: {10}(-272,132)(-272,160){11}
//: {12}(-118,132)(-118,184){13}
//: {14}(86,132)(86,181){15}
//: {16}(243,132)(243,185){17}
wire [3:0] w3;    //: /sn:0 {0}(-599,629)(-599,575){1}
//: {2}(-599,574)(-599,501)(-600,501)(-600,364){3}
//: {4}(-600,363)(-600,130){5}
//: {6}(-600,129)(-600,19){7}
//: {8}(-600,18)(-600,2){9}
wire w66;    //: /sn:0 /dp:1 {0}(79,284)(79,378)(37,378)(37,460){1}
wire w37;    //: /sn:0 {0}(157,420)(157,450)(58,450)(58,460){1}
wire w34;    //: /sn:0 {0}(-1,422)(-1,451)(-108,451)(-108,461){1}
wire w87;    //: /sn:0 /dp:1 {0}(-143,688)(-143,676)(-72,676)(-72,663){1}
wire w76;    //: /sn:0 {0}(-115,503)(-115,617)(8,617)(8,686){1}
wire w21;    //: /sn:0 {0}(-237,542)(-237,645){1}
wire w54;    //: /sn:0 {0}(259,575)(93,575){1}
//: {2}(89,575)(-64,575){3}
//: {4}(-68,575)(-227,575){5}
//: {6}(-231,575)(-423,575){7}
//: {8}(-427,575)(-595,575){9}
//: {10}(-425,577)(-425,611)(-428,611)(-428,638){11}
//: {12}(-229,577)(-229,615)(-232,615)(-232,645){13}
//: {14}(-66,577)(-66,613)(-69,613)(-69,642){15}
//: {16}(91,577)(91,610)(88,610)(88,636){17}
wire w31;    //: /sn:0 {0}(-162,423)(-162,453)(-266,453)(-266,463){1}
wire w28;    //: /sn:0 {0}(-314,405)(-314,442)(-436,442)(-436,465){1}
wire w41;    //: /sn:0 {0}(173,261)(140,261)(140,262)(99,262){1}
wire w20;    //: /sn:0 {0}(-76,541)(-76,632)(-74,632)(-74,642){1}
wire w36;    //: /sn:0 {0}(155,399)(155,348)(154,348)(154,340){1}
wire w1;    //: /sn:0 {0}(279,46)(279,54)(281,54)(281,64){1}
wire w25;    //: /sn:0 {0}(240,206)(240,224)(210,224)(210,234){1}
wire w74;    //: /sn:0 /dp:1 {0}(-95,481)(-71,481)(-71,487)(21,487){1}
wire w65;    //: /sn:0 {0}(57,264)(-68,264){1}
wire w92;    //: /sn:0 /dp:1 {0}(-320,686)(-320,676)(-235,676)(-235,666){1}
wire w91;    //: /sn:0 /dp:1 {0}(-150,730)(-150,806)(429,806){1}
wire w18;    //: /sn:0 {0}(-3,340)(-3,401){1}
wire w8;    //: /sn:0 {0}(-311,258)(-311,228)(-275,228)(-275,181){1}
wire w101;    //: /sn:0 /dp:1 {0}(-505,729)(-505,786)(429,786){1}
wire w71;    //: /sn:0 {0}(-88,286)(-88,423)(-124,423)(-124,461){1}
wire w30;    //: /sn:0 /dp:1 {0}(-164,402)(-164,348)(-165,348)(-165,340){1}
wire w17;    //: /sn:0 {0}(83,541)(83,636){1}
wire w22;    //: /sn:0 {0}(83,202)(83,232)(86,232)(86,242){1}
wire w84;    //: /sn:0 {0}(-423,485)(-295,485){1}
wire w59;    //: /sn:0 {0}(29,686)(29,670)(85,670)(85,657){1}
wire w85;    //: /sn:0 {0}(-465,487)(-485,487)(-485,649)(-514,649)(-514,687){1}
wire w57;    //: /sn:0 {0}(-301,309)(-301,450)(-282,450)(-282,463){1}
wire w12;    //: /sn:0 {0}(81,101)(81,181){1}
wire w11;    //: /sn:0 {0}(238,101)(238,185){1}
wire w2;    //: /sn:0 {0}(-165,80)(-165,232)(-97,232)(-97,244){1}
wire w70;    //: /sn:0 /dp:1 {0}(-110,266)(-223,266)(-223,246)(-290,246)(-290,258){1}
wire w10;    //: /sn:0 {0}(127,81)(127,224)(189,224)(189,234){1}
wire w94;    //: /sn:0 {0}(-307,706)(-182,706)(-182,710)(-172,710){1}
wire w27;    //: /sn:0 {0}(-316,384)(-316,358)(-319,358)(-319,340){1}
wire w13;    //: /sn:0 {0}(283,85)(283,846)(429,846){1}
wire w86;    //: /sn:0 {0}(-443,507)(-443,676)(-336,676)(-336,686){1}
wire w48;    //: /sn:0 {0}(47,511)(47,826)(429,826){1}
wire w52;    //: /sn:0 {0}(387,364)(162,364){1}
//: {2}(158,364)(3,364){3}
//: {4}(-1,364)(-158,364){5}
//: {6}(-162,364)(-309,364){7}
//: {8}(-311,362)(-311,384){9}
//: {10}(-313,364)(-596,364){11}
//: {12}(-160,366)(-160,376)(-159,376)(-159,402){13}
//: {14}(1,366)(1,376)(2,376)(2,401){15}
//: {16}(160,366)(160,399){17}
wire [3:0] w5;    //: /sn:0 {0}(340,97)(238,97){1}
//: {2}(237,97)(81,97){3}
//: {4}(80,97)(-123,97){5}
//: {6}(-124,97)(-279,97){7}
//: {8}(-280,97)(-499,97){9}
//: {10}(-501,95)(-501,44){11}
//: {12}(-499,42)(-171,42){13}
//: {14}(-170,42)(-91,42){15}
//: {16}(-90,42)(119,42){17}
//: {18}(120,42)(278,42){19}
//: {20}(279,42)(384,42){21}
//: {22}(-501,40)(-501,2){23}
//: {24}(-501,99)(-501,334){25}
//: {26}(-499,336)(-402,336)(-402,336)(-320,336){27}
//: {28}(-319,336)(-166,336){29}
//: {30}(-165,336)(-4,336){31}
//: {32}(-3,336)(153,336){33}
//: {34}(154,336)(223,336){35}
//: {36}(-501,338)(-501,536){37}
//: {38}(-499,538)(-431,538){39}
//: {40}(-430,538)(-238,538){41}
//: {42}(-237,538)(-162,538)(-162,537)(-77,537){43}
//: {44}(-76,537)(82,537){45}
//: {46}(83,537)(188,537){47}
//: {48}(-501,540)(-501,605){49}
wire w79;    //: /sn:0 {0}(-253,483)(-137,483){1}
wire w42;    //: /sn:0 {0}(200,285)(200,836)(429,836){1}
wire w50;    //: /sn:0 {0}(-167,59)(-167,54)(-170,54)(-170,46){1}
wire w9;    //: /sn:0 {0}(120,46)(120,54)(125,54)(125,60){1}
wire w26;    //: /sn:0 /dp:1 {0}(-121,205)(-121,225)(-81,225)(-81,244){1}
//: enddecls

  SHA g61 (.A(w70), .B(w8), .C(w56), .S(w57));   //: @(-326, 259) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  and g8 (.I0(w0), .I1(w12), .Z(w22));   //: @(83,192) /sn:0 /R:3 /w:[ 15 1 0 ]
  and g4 (.I0(w4), .I1(w9), .Z(w10));   //: @(127,71) /sn:0 /R:3 /w:[ 11 1 0 ]
  concat g58 (.I0(w13), .I1(w42), .I2(w48), .I3(w61), .I4(w91), .I5(w96), .I6(w101), .I7(w38), .Z(w19));   //: @(434,811) /sn:0 /w:[ 1 1 1 1 1 1 1 0 1 ] /dr:0
  tran g55(.Z(w20), .I(w5[1]));   //: @(-76,535) /sn:0 /R:1 /w:[ 0 43 44 ] /ss:1
  tran g51(.Z(w30), .I(w5[2]));   //: @(-165,334) /sn:0 /R:1 /w:[ 1 29 30 ] /ss:1
  //: joint g37 (w54) @(-229, 575) /w:[ 5 -1 6 12 ]
  //: joint g34 (w52) @(-311, 364) /w:[ 7 8 10 -1 ]
  and g13 (.I0(w52), .I1(w36), .Z(w37));   //: @(157,410) /sn:0 /R:3 /w:[ 17 0 0 ]
  and g3 (.I0(w4), .I1(w6), .Z(w7));   //: @(-85,72) /sn:0 /R:3 /w:[ 0 1 0 ]
  SFA g65 (.B(w71), .A(w34), .Ci(w74), .Co(w79), .S(w76));   //: @(-136, 462) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  //: dip g2 (w5) @(-501,-8) /sn:0 /w:[ 23 ] /st:2
  SHA g59 (.A(w25), .B(w10), .C(w41), .S(w42));   //: @(174, 235) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: dip g1 (w3) @(-600,-8) /sn:0 /w:[ 9 ] /st:8
  SFA g64 (.B(w2), .A(w26), .Ci(w65), .Co(w70), .S(w71));   //: @(-109, 245) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g16 (.I0(w54), .I1(w20), .Z(w87));   //: @(-72,653) /sn:0 /R:3 /w:[ 15 1 1 ]
  and g11 (.I0(w52), .I1(w30), .Z(w31));   //: @(-162,413) /sn:0 /R:3 /w:[ 13 0 0 ]
  tran g50(.Z(w18), .I(w5[1]));   //: @(-3,334) /sn:0 /R:1 /w:[ 0 31 32 ] /ss:1
  //: joint g28 (w0) @(-272, 130) /w:[ 7 -1 8 10 ]
  and g10 (.I0(w52), .I1(w27), .Z(w28));   //: @(-314,395) /sn:0 /R:3 /w:[ 9 0 0 ]
  //: joint g32 (w52) @(1, 364) /w:[ 3 -1 4 14 ]
  //: joint g27 (w0) @(243, 130) /w:[ 1 -1 2 16 ]
  //: joint g19 (w4) @(287, 19) /w:[ 6 -1 5 8 ]
  SFA g69 (.B(w86), .A(w92), .Ci(w94), .Co(w99), .S(w96));   //: @(-348, 687) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g38 (w54) @(-425, 575) /w:[ 7 -1 8 10 ]
  and g6 (.I0(w0), .I1(w15), .Z(w8));   //: @(-275,171) /sn:0 /R:3 /w:[ 11 1 1 ]
  //: joint g57 (w5) @(-501, 538) /w:[ 38 37 -1 48 ]
  tran g53(.Z(w51), .I(w5[3]));   //: @(-430,536) /sn:0 /R:1 /w:[ 0 39 40 ] /ss:1
  and g9 (.I0(w0), .I1(w11), .Z(w25));   //: @(240,196) /sn:0 /R:3 /w:[ 17 1 0 ]
  and g7 (.I0(w0), .I1(w14), .Z(w26));   //: @(-121,195) /sn:0 /R:3 /w:[ 13 1 0 ]
  led g71 (.I(w19));   //: @(536,74) /sn:0 /w:[ 0 ] /type:3
  //: joint g31 (w52) @(160, 364) /w:[ 1 -1 2 16 ]
  //: joint g20 (w4) @(130, 19) /w:[ 4 -1 3 10 ]
  and g15 (.I0(w54), .I1(w21), .Z(w92));   //: @(-235,656) /sn:0 /R:3 /w:[ 13 1 1 ]
  SFA g68 (.B(w16), .A(w87), .Ci(w89), .Co(w94), .S(w91));   //: @(-171, 689) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  SFA g67 (.B(w56), .A(w28), .Ci(w84), .Co(w85), .S(w86));   //: @(-464, 466) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  tran g39(.Z(w50), .I(w5[3]));   //: @(-170,40) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  tran g48(.Z(w27), .I(w5[3]));   //: @(-319,334) /sn:0 /R:1 /w:[ 1 27 28 ] /ss:1
  //: joint g43 (w5) @(-501, 97) /w:[ 9 10 -1 24 ]
  SHA g62 (.A(w59), .B(w76), .C(w89), .S(w61));   //: @(-7, 687) /sz:(47, 49) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<1 Bo0<0 ]
  //: joint g29 (w0) @(-118, 130) /w:[ 5 -1 6 12 ]
  tran g25(.Z(w54), .I(w3[3]));   //: @(-601,575) /sn:0 /R:2 /w:[ 9 1 2 ] /ss:1
  and g17 (.I0(w54), .I1(w17), .Z(w59));   //: @(85,647) /sn:0 /R:3 /w:[ 17 1 1 ]
  SFA g63 (.B(w7), .A(w22), .Ci(w41), .Co(w65), .S(w66));   //: @(58, 243) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g52 (w5) @(-501, 336) /w:[ 26 25 -1 36 ]
  tran g42(.Z(w1), .I(w5[0]));   //: @(279,40) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  tran g56(.Z(w21), .I(w5[2]));   //: @(-237,536) /sn:0 /R:1 /w:[ 0 41 42 ] /ss:1
  and g14 (.I0(w54), .I1(w51), .Z(w97));   //: @(-431,649) /sn:0 /R:3 /w:[ 11 1 1 ]
  and g5 (.I0(w4), .I1(w1), .Z(w13));   //: @(283,75) /sn:0 /R:3 /w:[ 9 1 0 ]
  tran g47(.Z(w15), .I(w5[3]));   //: @(-279,95) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  tran g44(.Z(w11), .I(w5[0]));   //: @(238,95) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g36 (w54) @(-66, 575) /w:[ 3 -1 4 14 ]
  //: joint g24 (w4) @(-162, 19) /w:[ 13 -1 14 16 ]
  tran g21(.Z(w0), .I(w3[1]));   //: @(-602,130) /sn:0 /R:2 /w:[ 9 5 6 ] /ss:1
  tran g41(.Z(w9), .I(w5[1]));   //: @(120,40) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  tran g23(.Z(w52), .I(w3[2]));   //: @(-602,364) /sn:0 /R:2 /w:[ 11 3 4 ] /ss:1
  SHA g60 (.A(w37), .B(w66), .C(w74), .S(w48));   //: @(22, 461) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  tran g54(.Z(w17), .I(w5[0]));   //: @(83,535) /sn:0 /R:1 /w:[ 0 45 46 ] /ss:1
  tran g40(.Z(w6), .I(w5[2]));   //: @(-90,40) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  SFA g70 (.B(w85), .A(w97), .Ci(w99), .Co(w38), .S(w101));   //: @(-526, 688) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  tran g46(.Z(w14), .I(w5[2]));   //: @(-123,95) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g45(.Z(w12), .I(w5[1]));   //: @(81,95) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: joint g35 (w54) @(91, 575) /w:[ 1 -1 2 16 ]
  //: joint g26 (w5) @(-501, 42) /w:[ 12 22 -1 11 ]
  //: joint g22 (w4) @(-82, 19) /w:[ 2 -1 12 1 ]
  and g0 (.I0(w4), .I1(w50), .Z(w2));   //: @(-165,70) /sn:0 /R:3 /w:[ 17 0 0 ]
  SFA g66 (.B(w57), .A(w31), .Ci(w79), .Co(w84), .S(w16));   //: @(-294, 464) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  tran g18(.Z(w4), .I(w3[0]));   //: @(-602,19) /sn:0 /R:2 /w:[ 15 7 8 ] /ss:1
  and g12 (.I0(w52), .I1(w18), .Z(w34));   //: @(-1,412) /sn:0 /R:3 /w:[ 15 1 0 ]
  //: joint g33 (w52) @(-160, 364) /w:[ 5 -1 6 12 ]
  //: joint g30 (w0) @(86, 130) /w:[ 3 -1 4 14 ]
  tran g49(.Z(w36), .I(w5[0]));   //: @(154,334) /sn:0 /R:1 /w:[ 1 33 34 ] /ss:1

endmodule

module SHA(S, B, A, C);
//: interface  /sz:(47, 49) /bd:[ Ti0>B(15/47) Ti1>A(36/47) Lo0<C(26/49) Bo0<S(26/47) ]
input B;    //: /sn:0 {0}(97,314)(228,314)(228,308){1}
//: {2}(230,306)(240,306)(240,311)(296,311){3}
//: {4}(228,304)(228,252)(296,252){5}
input A;    //: /sn:0 {0}(115,248)(244,248){1}
//: {2}(248,248)(288,248)(288,247)(296,247){3}
//: {4}(246,250)(246,306)(296,306){5}
output C;    //: /sn:0 {0}(469,310)(327,310)(327,309)(317,309){1}
output S;    //: /sn:0 /dp:1 {0}(317,250)(459,250)(459,253)(469,253){1}
//: enddecls

  //: output g4 (S) @(466,253) /sn:0 /w:[ 1 ]
  //: input g3 (B) @(95,314) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(113,248) /sn:0 /w:[ 0 ]
  and g1 (.I0(A), .I1(B), .Z(C));   //: @(307,309) /sn:0 /w:[ 5 3 1 ]
  //: joint g6 (B) @(228, 306) /w:[ 2 4 -1 1 ]
  //: joint g7 (A) @(246, 248) /w:[ 2 -1 1 4 ]
  //: output g5 (C) @(466,310) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(S));   //: @(307,250) /sn:0 /w:[ 3 5 0 ]

endmodule
