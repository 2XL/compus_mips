//: version "1.8.7"

module main;    //: root_module
wire w32;    //: /sn:0 /dp:1 {0}(416,216)(416,267)(954,267){1}
wire w6;    //: /sn:0 {0}(954,307)(750,307)(750,216){1}
wire w7;    //: /sn:0 {0}(769,192)(811,192){1}
wire w14;    //: /sn:0 {0}(507,128)(507,136)(504,136)(504,174){1}
wire w16;    //: /sn:0 {0}(922,128)(922,174){1}
wire [7:0] w4;    //: /sn:0 /dp:9 {0}(72,110)(72,124)(337,124){1}
//: {2}(338,124)(423,124){3}
//: {4}(424,124)(506,124){5}
//: {6}(507,124)(587,124){7}
//: {8}(588,124)(670,124){9}
//: {10}(671,124)(753,124){11}
//: {12}(754,124)(837,124){13}
//: {14}(838,124)(921,124){15}
//: {16}(922,124)(1060,124){17}
wire w19;    //: /sn:0 {0}(352,192)(393,192){1}
wire w15;    //: /sn:0 {0}(838,128)(838,174){1}
wire w38;    //: /sn:0 {0}(572,68)(572,76)(577,76)(577,174){1}
wire w3;    //: /sn:0 {0}(671,128)(671,174){1}
wire w0;    //: /sn:0 {0}(660,68)(660,174){1}
wire w34;    //: /sn:0 {0}(338,128)(338,136)(337,136)(337,174){1}
wire [8:0] w21;    //: /sn:0 /dp:1 {0}(960,287)(1053,287){1}
wire w31;    //: /sn:0 {0}(409,68)(409,174){1}
wire w28;    //: /sn:0 {0}(519,192)(561,192){1}
wire [7:0] w24;    //: /sn:0 /dp:17 {0}(1053,64)(911,64){1}
//: {2}(910,64)(827,64){3}
//: {4}(826,64)(743,64){5}
//: {6}(742,64)(660,64){7}
//: {8}(659,64)(572,64){9}
//: {10}(571,64)(489,64){11}
//: {12}(488,64)(409,64){13}
//: {14}(408,64)(325,64){15}
//: {16}(324,64)(72,64)(72,59){17}
wire w23;    //: /sn:0 /dp:1 {0}(333,216)(333,257)(954,257){1}
wire w20;    //: /sn:0 /dp:1 {0}(954,317)(834,317)(834,216){1}
wire w1;    //: /sn:0 {0}(743,68)(743,174){1}
wire w25;    //: /sn:0 {0}(489,68)(489,76)(493,76)(493,174){1}
wire w35;    //: /sn:0 {0}(603,192)(644,192){1}
wire w18;    //: /sn:0 /dp:1 {0}(954,327)(918,327)(918,216){1}
wire w8;    //: /sn:0 {0}(686,192)(727,192){1}
wire w30;    //: /sn:0 /dp:1 {0}(584,216)(584,287)(954,287){1}
wire w17;    //: /sn:0 {0}(435,192)(477,192){1}
wire w22;    //: /sn:0 {0}(954,297)(667,297)(667,216){1}
wire w2;    //: /sn:0 {0}(325,68)(325,76)(326,76)(326,174){1}
wire w11;    //: /sn:0 {0}(754,128)(754,174){1}
wire w12;    //: /sn:0 {0}(911,68)(911,174){1}
wire w10;    //: /sn:0 {0}(91,180)(91,192)(211,192){1}
//: {2}(215,192)(310,192){3}
//: {4}(213,194)(213,247)(954,247){5}
wire w13;    //: /sn:0 {0}(853,192)(895,192){1}
wire w33;    //: /sn:0 {0}(424,128)(424,136)(420,136)(420,174){1}
wire w5;    //: /sn:0 {0}(976,192)(937,192){1}
wire w29;    //: /sn:0 /dp:1 {0}(500,216)(500,277)(954,277){1}
wire w9;    //: /sn:0 {0}(827,68)(827,174){1}
wire w26;    //: /sn:0 {0}(588,128)(588,174){1}
//: enddecls

  led g8 (.I(w10));   //: @(91,173) /sn:0 /w:[ 0 ] /type:0
  SFA g4 (.B(w11), .A(w1), .Ci(w7), .Co(w8), .S(w6));   //: @(728, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  tran g13(.Z(w9), .I(w24[1]));   //: @(827,62) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  tran g3(.Z(w0), .I(w24[3]));   //: @(660,62) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  led g2 (.I(w21));   //: @(1060,287) /sn:0 /R:3 /w:[ 1 ] /type:3
  //: dip g1 (w24) @(72,49) /sn:0 /w:[ 17 ] /st:9
  tran g16(.Z(w16), .I(w4[0]));   //: @(922,122) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  tran g11(.Z(w1), .I(w24[2]));   //: @(743,62) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  tran g28(.Z(w14), .I(w4[5]));   //: @(507,122) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g10(.Z(w3), .I(w4[3]));   //: @(671,122) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  tran g27(.Z(w33), .I(w4[6]));   //: @(424,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g19(.Z(w25), .I(w24[5]));   //: @(489,62) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  SFA g6 (.B(w16), .A(w12), .Ci(w5), .Co(w13), .S(w18));   //: @(896, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  //: dip g9 (w4) @(72,100) /sn:0 /w:[ 0 ] /st:0
  concat g7 (.I0(w18), .I1(w20), .I2(w6), .I3(w22), .I4(w30), .I5(w29), .I6(w32), .I7(w23), .I8(w10), .Z(w21));   //: @(959,287) /sn:0 /w:[ 0 0 0 0 1 1 1 1 5 0 ] /dr:0
  SFA g20 (.B(w33), .A(w31), .Ci(w17), .Co(w19), .S(w32));   //: @(394, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  tran g15(.Z(w15), .I(w4[1]));   //: @(838,122) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  tran g29(.Z(w26), .I(w4[4]));   //: @(588,122) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g25(.Z(w2), .I(w24[7]));   //: @(325,62) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  //: switch g17 (w5) @(994,192) /sn:0 /R:2 /w:[ 0 ] /st:0
  tran g14(.Z(w12), .I(w24[0]));   //: @(911,62) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  SFA g5 (.B(w15), .A(w9), .Ci(w13), .Co(w7), .S(w20));   //: @(812, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  tran g24(.Z(w31), .I(w24[6]));   //: @(409,62) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  SFA g21 (.B(w26), .A(w38), .Ci(w35), .Co(w28), .S(w30));   //: @(562, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  SFA g23 (.B(w34), .A(w2), .Ci(w19), .Co(w10), .S(w23));   //: @(311, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<3 Bo0<0 ]
  tran g26(.Z(w34), .I(w4[7]));   //: @(338,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  SFA g22 (.B(w14), .A(w25), .Ci(w28), .Co(w17), .S(w29));   //: @(478, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  SFA g0 (.B(w3), .A(w0), .Ci(w8), .Co(w35), .S(w22));   //: @(645, 175) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]
  tran g18(.Z(w38), .I(w24[4]));   //: @(572,62) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  tran g12(.Z(w11), .I(w4[2]));   //: @(754,122) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  //: joint g30 (w10) @(213, 192) /w:[ 2 -1 1 4 ]

endmodule

module SFA(S, Ci, B, A, Co);
//: interface  /sz:(40, 40) /bd:[ Ti0>A(15/40) Ti1>B(26/40) Ri0>Ci(17/40) Lo0<Co(17/40) Bo0<S(22/40) ]
input B;    //: /sn:0 {0}(66,121)(105,121){1}
//: {2}(109,121)(149,121)(149,103)(157,103){3}
//: {4}(107,123)(107,193)(163,193){5}
input A;    //: /sn:0 /dp:1 {0}(157,98)(99,98)(99,102){1}
//: {2}(97,104)(65,104){3}
//: {4}(99,106)(99,188)(163,188){5}
output Co;    //: /sn:0 {0}(288,178)(249,178){1}
input Ci;    //: /sn:0 {0}(67,141)(132,141){1}
//: {2}(136,141)(212,141)(212,127)(220,127){3}
//: {4}(134,143)(134,162)(164,162){5}
output S;    //: /sn:0 {0}(286,125)(241,125){1}
wire w8;    //: /sn:0 {0}(184,191)(218,191)(218,180)(228,180){1}
wire w2;    //: /sn:0 {0}(178,101)(190,101){1}
//: {2}(194,101)(210,101)(210,122)(220,122){3}
//: {4}(192,103)(192,132)(155,132)(155,167)(164,167){5}
wire w5;    //: /sn:0 {0}(185,165)(218,165)(218,175)(228,175){1}
//: enddecls

  //: joint g8 (A) @(99, 104) /w:[ -1 1 2 4 ]
  and g4 (.I0(Ci), .I1(w2), .Z(w5));   //: @(175,165) /sn:0 /w:[ 5 5 0 ]
  //: output g13 (S) @(283,125) /sn:0 /w:[ 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(168,101) /sn:0 /w:[ 0 3 0 ]
  //: input g2 (Ci) @(65,141) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(64,121) /sn:0 /w:[ 0 ]
  //: joint g11 (w2) @(192, 101) /w:[ 2 -1 1 4 ]
  //: joint g10 (Ci) @(134, 141) /w:[ 2 -1 1 4 ]
  or g6 (.I0(w5), .I1(w8), .Z(Co));   //: @(239,178) /sn:0 /w:[ 1 1 1 ]
  //: joint g9 (B) @(107, 121) /w:[ 2 -1 1 4 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(S));   //: @(231,125) /sn:0 /w:[ 3 3 1 ]
  and g5 (.I0(A), .I1(B), .Z(w8));   //: @(174,191) /sn:0 /w:[ 5 5 0 ]
  //: input g0 (A) @(63,104) /sn:0 /w:[ 3 ]
  //: output g12 (Co) @(285,178) /sn:0 /w:[ 0 ]

endmodule
