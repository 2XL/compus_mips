//: version "1.8.7"

module main;    //: root_module
wire w96;    //: /sn:0 {0}(893,402)(893,410)(908,410)(908,270)(934,270)(934,294){1}
wire w93;    //: /sn:0 {0}(912,166)(912,175)(1045,175)(1045,209){1}
wire w7;    //: /sn:0 {0}(918,312)(879,312)(879,433)(859,433){1}
wire w45;    //: /sn:0 {0}(242,545)(232,545)(232,617)(1226,617){1}
wire w99;    //: /sn:0 {0}(293,401)(293,426)(370,426)(370,436){1}
wire w60;    //: /sn:0 /dp:1 {0}(859,210)(859,172)(695,172)(695,165){1}
wire w46;    //: /sn:0 {0}(265,569)(265,627)(1226,627){1}
wire [3:0] w56;    //: /sn:0 {0}(115,-41)(170,-41){1}
//: {2}(171,-41)(199,-41){3}
//: {4}(200,-41)(227,-41){5}
//: {6}(228,-41)(260,-41){7}
//: {8}(261,-41)(1224,-41){9}
wire w16;    //: /sn:0 /dp:1 {0}(648,259)(648,282)(709,282)(709,298){1}
wire w81;    //: /sn:0 {0}(446,488)(446,498)(431,498)(431,425)(381,425)(381,436){1}
wire w19;    //: /sn:0 {0}(1226,667)(941,667)(941,336){1}
wire w15;    //: /sn:0 /dp:1 {0}(622,233)(593,233)(593,323)(540,323){1}
wire w69;    //: /sn:0 {0}(413,293)(413,303)(428,303)(428,291)(514,291)(514,305){1}
wire w51;    //: /sn:0 {0}(492,574)(492,637)(1226,637){1}
wire w3;    //: /sn:0 /dp:1 {0}(1029,236)(1006,236)(1006,312)(960,312){1}
wire w66;    //: /sn:0 {0}(759,293)(759,303)(774,303)(774,164)(838,164)(838,210){1}
wire w64;    //: /sn:0 {0}(762,272)(762,60)(761,60)(761,61){1}
//: {2}(763,63)(978,63){3}
//: {4}(982,63)(1223,63){5}
//: {6}(980,65)(980,75)(981,75)(981,270){7}
//: {8}(759,63)(563,63){9}
//: {10}(559,63)(442,63){11}
//: {12}(438,63)(131,63)(131,41){13}
//: {14}(440,65)(440,75)(416,75)(416,272){15}
//: {16}(561,65)(561,272){17}
wire w63;    //: /sn:0 {0}(558,293)(558,294)(580,294)(580,182)(659,182)(659,205){1}
wire w102;    //: /sn:0 {0}(487,380)(487,385)(549,385)(549,263)(525,263)(525,305){1}
wire w87;    //: /sn:0 {0}(1124,170)(1124,687)(1226,687){1}
wire w21;    //: /sn:0 {0}(716,340)(716,405)(833,405)(833,415){1}
wire w54;    //: /sn:0 /dp:1 {0}(665,558)(511,558)(511,522)(496,522)(496,532){1}
wire w90;    //: /sn:0 {0}(571,166)(571,167)(593,167)(593,155)(638,155)(638,205){1}
wire w31;    //: /sn:0 {0}(840,457)(840,657)(1226,657){1}
wire w28;    //: /sn:0 {0}(844,415)(844,391)(803,391)(803,515)(788,515)(788,505){1}
wire w20;    //: /sn:0 {0}(693,316)(594,316)(594,429)(584,429){1}
wire w36;    //: /sn:0 {0}(566,453)(566,521)(681,521)(681,531){1}
wire w41;    //: /sn:0 {0}(377,478)(377,522)(485,522)(485,532){1}
wire w25;    //: /sn:0 {0}(498,323)(406,323)(406,454)(396,454){1}
wire w65;    //: /sn:0 {0}(757,272)(757,-6)(764,-6)(764,-14){1}
//: {2}(766,-16)(908,-16){3}
//: {4}(912,-16)(1224,-16){5}
//: {6}(910,-14)(910,-4)(915,-4)(915,145){7}
//: {8}(762,-16)(679,-16){9}
//: {10}(675,-16)(617,-16){11}
//: {12}(613,-16)(228,-16)(228,-37){13}
//: {14}(615,-14)(615,-4)(605,-4)(605,486){15}
//: {16}(677,-14)(677,186)(670,186)(670,350){17}
wire w103;    //: /sn:0 {0}(675,350)(675,193)(691,193)(691,174)(655,174)(655,77){1}
//: {2}(657,75)(892,75){3}
//: {4}(896,75)(1136,75){5}
//: {6}(894,77)(894,87)(896,87)(896,381){7}
//: {8}(653,75)(494,75){9}
//: {10}(490,75)(307,75){11}
//: {12}(303,75)(101,75)(101,41){13}
//: {14}(305,77)(305,87)(296,87)(296,380){15}
//: {16}(492,77)(492,214)(490,214)(490,359){17}
wire w35;    //: /sn:0 {0}(542,429)(523,429)(523,550)(511,550){1}
wire w40;    //: /sn:0 {0}(354,454)(294,454)(294,545)(284,545){1}
wire w71;    //: /sn:0 {0}(976,270)(976,-24)(979,-24)(979,-26){1}
//: {2}(981,-28)(1125,-28){3}
//: {4}(1129,-28)(1225,-28){5}
//: {6}(1127,-26)(1127,149){7}
//: {8}(977,-28)(877,-28){9}
//: {10}(873,-28)(795,-28){11}
//: {12}(791,-28)(261,-28)(261,-37){13}
//: {14}(793,-26)(793,-16)(786,-16)(786,484){15}
//: {16}(875,-26)(875,-16)(891,-16)(891,381){17}
wire w68;    //: /sn:0 {0}(171,-37)(171,7)(211,7){1}
//: {2}(215,7)(288,7){3}
//: {4}(292,7)(420,7){5}
//: {6}(424,7)(568,7){7}
//: {8}(572,7)(1224,7){9}
//: {10}(570,9)(570,19)(569,19)(569,145){11}
//: {12}(422,9)(422,19)(411,19)(411,272){13}
//: {14}(290,9)(290,19)(291,19)(291,380){15}
//: {16}(213,9)(213,19)(216,19)(216,480){17}
wire w30;    //: /sn:0 {0}(817,433)(702,433)(702,531){1}
wire w84;    //: /sn:0 {0}(218,501)(218,517)(258,517)(258,527){1}
wire w62;    //: /sn:0 {0}(556,272)(556,1)(529,1)(529,-2){1}
//: {2}(531,-4)(692,-4){3}
//: {4}(696,-4)(1226,-4){5}
//: {6}(694,-2)(694,8)(693,8)(693,144){7}
//: {8}(527,-4)(486,-4){9}
//: {10}(482,-4)(461,-4){11}
//: {12}(459,-6)(459,-21)(444,-21)(444,467){13}
//: {14}(457,-4)(200,-4)(200,-37){15}
//: {16}(484,-2)(484,162)(485,162)(485,359){17}
wire w2;    //: /sn:0 {0}(1055,260)(1055,677)(1226,677){1}
wire w11;    //: /sn:0 /dp:1 {0}(822,237)(779,237)(779,316)(735,316){1}
wire w12;    //: /sn:0 /dp:1 {0}(848,261)(848,284)(945,284)(945,294){1}
wire [3:0] w57;    //: /sn:0 {0}(6,37)(75,37){1}
//: {2}(76,37)(100,37){3}
//: {4}(101,37)(130,37){5}
//: {6}(131,37)(150,37){7}
//: {8}(151,37)(1137,37){9}
wire w110;    //: /sn:0 {0}(1133,90)(797,90){1}
//: {2}(793,90)(610,90){3}
//: {4}(606,90)(453,90){5}
//: {6}(451,88)(451,73)(449,73)(449,467){7}
//: {8}(449,90)(224,90){9}
//: {10}(220,90)(76,90)(76,41){11}
//: {12}(222,92)(222,102)(221,102)(221,480){13}
//: {14}(608,92)(608,102)(610,102)(610,486){15}
//: {16}(795,92)(795,102)(791,102)(791,484){17}
wire w105;    //: /sn:0 {0}(672,371)(672,381)(687,381)(687,240)(720,240)(720,298){1}
wire w78;    //: /sn:0 {0}(607,507)(607,517)(643,517)(643,403)(569,403)(569,411){1}
wire w72;    //: /sn:0 {0}(978,291)(978,301)(993,301)(993,142)(1066,142)(1066,209){1}
wire w52;    //: /sn:0 {0}(698,144)(698,40)(705,40)(705,50){1}
//: {2}(707,52)(908,52){3}
//: {4}(912,52)(1120,52){5}
//: {6}(1124,52)(1227,52){7}
//: {8}(1122,54)(1122,149){9}
//: {10}(910,54)(910,145){11}
//: {12}(703,52)(581,52){13}
//: {14}(577,52)(151,52)(151,41){15}
//: {16}(579,54)(579,64)(574,64)(574,145){17}
wire [7:0] w29;    //: /sn:0 /dp:1 {0}(1278,646)(1278,652)(1232,652){1}
wire w50;    //: /sn:0 {0}(469,550)(284,550)(284,517)(269,517)(269,527){1}
wire w26;    //: /sn:0 {0}(521,347)(521,401)(558,401)(558,411){1}
wire w55;    //: /sn:0 /dp:1 {0}(691,582)(691,647)(1226,647){1}
//: enddecls

  //: joint g61 (w103) @(492, 75) /w:[ 9 -1 10 16 ]
  SFA g4 (.B(w105), .A(w16), .Ci(w11), .Co(w20), .S(w21));   //: @(694, 299) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  SFA g8 (.B(w81), .A(w99), .Ci(w25), .Co(w40), .S(w41));   //: @(355, 437) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g58 (w103) @(655, 75) /w:[ 2 -1 8 1 ]
  //: joint g55 (w64) @(440, 63) /w:[ 11 -1 12 14 ]
  //: joint g51 (w65) @(764, -16) /w:[ 2 -1 8 1 ]
  tran g37(.Z(w110), .I(w57[3]));   //: @(76,35) /sn:0 /R:1 /w:[ 11 1 2 ] /ss:1
  tran g34(.Z(w62), .I(w56[2]));   //: @(200,-43) /sn:0 /R:1 /w:[ 15 3 4 ] /ss:1
  //: dip g13 (w57) @(-32,37) /sn:0 /R:1 /w:[ 0 ] /st:2
  SHA g3 (.B(w90), .A(w63), .C(w15), .S(w16));   //: @(623, 206) /sz:(47, 52) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g65 (w110) @(608, 90) /w:[ 3 -1 4 14 ]
  SHA g2 (.B(w66), .A(w60), .C(w11), .S(w12));   //: @(823, 211) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  //: joint g59 (w65) @(677, -16) /w:[ 9 -1 10 16 ]
  SFA g1 (.B(w12), .A(w96), .Ci(w3), .Co(w7), .S(w19));   //: @(919, 295) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g64 (w110) @(795, 90) /w:[ 1 -1 2 16 ]
  //: joint g16 (w71) @(1127, -28) /w:[ 4 -1 3 6 ]
  SHA g11 (.B(w36), .A(w30), .C(w54), .S(w55));   //: @(666, 532) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g50 (w64) @(761, 63) /w:[ 2 1 8 -1 ]
  and g28 (.I0(w52), .I1(w68), .Z(w90));   //: @(571,156) /sn:0 /R:3 /w:[ 17 11 0 ]
  SFA g10 (.B(w54), .A(w41), .Ci(w35), .Co(w50), .S(w51));   //: @(470, 533) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g32 (.I0(w103), .I1(w62), .Z(w102));   //: @(487,370) /sn:0 /R:3 /w:[ 17 17 0 ]
  and g27 (.I0(w71), .I1(w52), .Z(w87));   //: @(1124,160) /sn:0 /R:3 /w:[ 7 9 0 ]
  and g19 (.I0(w64), .I1(w62), .Z(w63));   //: @(558,283) /sn:0 /R:3 /w:[ 17 0 0 ]
  //: joint g69 (w65) @(615, -16) /w:[ 11 -1 12 14 ]
  //: joint g38 (w52) @(1122, 52) /w:[ 6 -1 5 8 ]
  SFA g6 (.B(w28), .A(w21), .Ci(w7), .Co(w30), .S(w31));   //: @(818, 416) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g57 (w71) @(875, -28) /w:[ 9 -1 10 16 ]
  //: joint g53 (w62) @(529, -4) /w:[ 2 -1 8 1 ]
  SFA g7 (.B(w78), .A(w26), .Ci(w20), .Co(w35), .S(w36));   //: @(543, 412) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  SFA g9 (.B(w50), .A(w84), .Ci(w40), .Co(w45), .S(w46));   //: @(243, 528) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g71 (w68) @(213, 7) /w:[ 2 -1 1 16 ]
  tran g15(.Z(w68), .I(w56[3]));   //: @(171,-43) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  and g31 (.I0(w103), .I1(w68), .Z(w99));   //: @(293,391) /sn:0 /R:3 /w:[ 15 15 0 ]
  and g20 (.I0(w64), .I1(w65), .Z(w66));   //: @(759,283) /sn:0 /R:3 /w:[ 0 0 0 ]
  //: joint g68 (w71) @(793, -28) /w:[ 11 -1 12 14 ]
  //: joint g67 (w110) @(222, 90) /w:[ 9 -1 10 12 ]
  tran g39(.Z(w103), .I(w57[2]));   //: @(101,35) /sn:0 /R:1 /w:[ 13 3 4 ] /ss:1
  //: joint g48 (w64) @(980, 63) /w:[ 4 -1 3 6 ]
  tran g43(.Z(w52), .I(w57[0]));   //: @(151,35) /sn:0 /R:1 /w:[ 15 7 8 ] /ss:1
  //: joint g62 (w68) @(290, 7) /w:[ 4 -1 3 14 ]
  and g29 (.I0(w65), .I1(w52), .Z(w93));   //: @(912,156) /sn:0 /R:3 /w:[ 7 11 0 ]
  and g25 (.I0(w110), .I1(w62), .Z(w81));   //: @(446,478) /sn:0 /R:3 /w:[ 7 13 0 ]
  led g17 (.I(w29));   //: @(1278,639) /sn:0 /w:[ 0 ] /type:2
  //: joint g63 (w103) @(305, 75) /w:[ 11 -1 12 14 ]
  //: joint g52 (w64) @(561, 63) /w:[ 9 -1 10 16 ]
  //: joint g42 (w52) @(910, 52) /w:[ 4 -1 3 10 ]
  //: joint g56 (w103) @(894, 75) /w:[ 4 -1 3 6 ]
  SFA g5 (.B(w102), .A(w69), .Ci(w15), .Co(w25), .S(w26));   //: @(499, 306) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  concat g14 (.I0(w87), .I1(w2), .I2(w19), .I3(w31), .I4(w55), .I5(w51), .I6(w46), .I7(w45), .Z(w29));   //: @(1231,652) /sn:0 /w:[ 1 1 0 1 1 1 1 1 1 ] /dr:0
  //: joint g47 (w52) @(579, 52) /w:[ 13 -1 14 16 ]
  //: joint g44 (w62) @(694, -4) /w:[ 4 -1 3 6 ]
  tran g36(.Z(w71), .I(w56[0]));   //: @(261,-43) /sn:0 /R:1 /w:[ 13 7 8 ] /ss:1
  and g24 (.I0(w110), .I1(w65), .Z(w78));   //: @(607,497) /sn:0 /R:3 /w:[ 15 15 0 ]
  and g21 (.I0(w64), .I1(w68), .Z(w69));   //: @(413,283) /sn:0 /R:3 /w:[ 15 13 0 ]
  tran g41(.Z(w64), .I(w57[1]));   //: @(131,35) /sn:0 /R:1 /w:[ 13 5 6 ] /ss:1
  and g23 (.I0(w110), .I1(w71), .Z(w28));   //: @(788,495) /sn:0 /R:3 /w:[ 17 15 1 ]
  //: joint g60 (w62) @(484, -4) /w:[ 9 -1 10 16 ]
  //: joint g54 (w68) @(422, 7) /w:[ 6 -1 5 12 ]
  //: joint g40 (w65) @(910, -16) /w:[ 4 -1 3 6 ]
  //: joint g70 (w62) @(459, -4) /w:[ 11 12 14 -1 ]
  //: joint g46 (w68) @(570, 7) /w:[ 8 -1 7 10 ]
  //: joint g45 (w52) @(705, 52) /w:[ 2 1 12 -1 ]
  tran g35(.Z(w65), .I(w56[1]));   //: @(228,-43) /sn:0 /R:1 /w:[ 13 5 6 ] /ss:1
  and g26 (.I0(w110), .I1(w68), .Z(w84));   //: @(218,491) /sn:0 /R:3 /w:[ 13 17 0 ]
  and g22 (.I0(w64), .I1(w71), .Z(w72));   //: @(978,281) /sn:0 /R:3 /w:[ 7 0 0 ]
  SHA g0 (.B(w93), .A(w72), .C(w3), .S(w2));   //: @(1030, 210) /sz:(47, 49) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g66 (w110) @(451, 90) /w:[ 5 6 8 -1 ]
  and g18 (.I0(w52), .I1(w62), .Z(w60));   //: @(695,155) /sn:0 /R:3 /w:[ 0 7 1 ]
  //: dip g12 (w56) @(77,-41) /sn:0 /R:1 /w:[ 0 ] /st:8
  and g33 (.I0(w103), .I1(w65), .Z(w105));   //: @(672,361) /sn:0 /R:3 /w:[ 0 17 0 ]
  and g30 (.I0(w103), .I1(w71), .Z(w96));   //: @(893,392) /sn:0 /R:3 /w:[ 7 17 0 ]
  //: joint g49 (w71) @(979, -28) /w:[ 2 -1 8 1 ]

endmodule

module SHA(S, B, A, C);
//: interface  /sz:(47, 49) /bd:[ Ti0>B(15/47) Ti1>A(36/47) Lo0<C(26/49) Bo0<S(25/47) ]
input B;    //: /sn:0 {0}(129,181)(260,181)(260,175){1}
//: {2}(262,173)(272,173)(272,178)(328,178){3}
//: {4}(260,171)(260,119)(328,119){5}
input A;    //: /sn:0 {0}(147,115)(276,115){1}
//: {2}(280,115)(320,115)(320,114)(328,114){3}
//: {4}(278,117)(278,173)(328,173){5}
output C;    //: /sn:0 {0}(501,177)(359,177)(359,176)(349,176){1}
output S;    //: /sn:0 {0}(349,117)(491,117)(491,120)(501,120){1}
//: enddecls

  //: output g4 (S) @(498,120) /sn:0 /w:[ 1 ]
  //: input g3 (B) @(127,181) /sn:0 /w:[ 0 ]
  //: input g2 (A) @(145,115) /sn:0 /w:[ 0 ]
  and g1 (.I0(A), .I1(B), .Z(C));   //: @(339,176) /sn:0 /w:[ 5 3 1 ]
  //: joint g6 (B) @(260, 173) /w:[ 2 4 -1 1 ]
  //: joint g7 (A) @(278, 115) /w:[ 2 -1 1 4 ]
  //: output g5 (C) @(498,177) /sn:0 /w:[ 0 ]
  xor g0 (.I0(A), .I1(B), .Z(S));   //: @(339,117) /sn:0 /w:[ 3 5 0 ]

endmodule
