//: version "1.8.7"

module main;    //: root_module
wire A;    //: /sn:0 /dp:1 {0}(-447,54)(-58,54)(-58,207)(-45,207)(-45,242)(178,242)(178,256){1}
wire G;    //: /sn:0 /dp:1 {0}(69,366)(33,366)(33,511)(195,511)(195,298){1}
wire [2:0] w28;    //: /sn:0 {0}(314,324)(314,537)(104,537)(104,356)(75,356){1}
wire P;    //: /sn:0 /dp:1 {0}(69,356)(-13,356)(-13,424)(186,424)(186,298){1}
wire C;    //: /sn:0 {0}(-446,188)(211,188)(211,246)(191,246)(191,256){1}
wire w29;    //: /sn:0 {0}(205,276)(241,276)(241,129)(-230,129)(-230,118)(-447,118){1}
wire S;    //: /sn:0 {0}(69,346)(38,346)(38,313)(176,313)(176,298){1}
//: enddecls

  //: switch g13 (C) @(-463,188) /sn:0 /w:[ 0 ] /st:0
  concat g11 (.I0(G), .I1(P), .I2(S), .Z(w28));   //: @(74,356) /sn:0 /w:[ 0 0 0 1 ] /dr:0
  led g10 (.I(w28));   //: @(314,317) /sn:0 /w:[ 0 ] /type:2
  //: switch g9 (A) @(-464,54) /sn:0 /w:[ 0 ] /st:0
  S_CLA g17 (.A(A), .B(C), .C(w29), .P(S), .G(P), .S(G));   //: @(164, 257) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]
  //: switch g12 (w29) @(-464,118) /sn:0 /w:[ 1 ] /st:0

endmodule

module S_CLA(G, S, P, A, B, C);
//: interface  /sz:(40, 40) /bd:[ Ti0>B(27/40) Ti1>A(14/40) Ri0>C(19/40) Bo0<S(31/40) Bo1<G(22/40) Bo2<P(12/40) ]
input B;    //: /sn:0 {0}(82,131)(125,131){1}
//: {2}(129,131)(152,131)(152,121)(226,121){3}
//: {4}(127,133)(127,152){5}
//: {6}(129,154)(340,154){7}
//: {8}(127,156)(127,192)(339,192){9}
input A;    //: /sn:0 {0}(81,107)(102,107){1}
//: {2}(106,107)(153,107)(153,116)(226,116){3}
//: {4}(104,109)(104,120)(117,120)(117,153){5}
//: {6}(119,155)(236,155)(236,159)(340,159){7}
//: {8}(117,157)(117,197)(339,197){9}
output G;    //: /sn:0 {0}(360,195)(448,195){1}
output P;    //: /sn:0 /dp:1 {0}(361,157)(448,157){1}
input C;    //: /sn:0 {0}(37,146)(270,146)(270,106)(338,106){1}
output S;    //: /sn:0 {0}(359,104)(448,104){1}
wire w3;    //: /sn:0 {0}(338,101)(299,101)(299,119)(247,119){1}
//: enddecls

  xor g34 (.I0(A), .I1(B), .Z(w3));   //: @(237,119) /sn:0 /w:[ 3 3 1 ]
  //: joint g28 (A) @(117, 155) /w:[ 6 5 -1 8 ]
  //: output g32 (G) @(445,195) /sn:0 /w:[ 1 ]
  xor g27 (.I0(w3), .I1(C), .Z(S));   //: @(349,104) /sn:0 /w:[ 0 1 0 ]
  //: output g31 (S) @(445,104) /sn:0 /w:[ 1 ]
  //: joint g29 (A) @(104, 107) /w:[ 2 -1 1 4 ]
  //: joint g25 (B) @(127, 154) /w:[ 6 5 -1 8 ]
  and g24 (.I0(B), .I1(A), .Z(G));   //: @(350,195) /sn:0 /w:[ 9 9 0 ]
  //: output g23 (P) @(445,157) /sn:0 /w:[ 1 ]
  //: joint g35 (B) @(127, 131) /w:[ 2 -1 1 4 ]
  or g26 (.I0(B), .I1(A), .Z(P));   //: @(351,157) /sn:0 /w:[ 7 7 0 ]
  //: input g22 (A) @(79,107) /sn:0 /w:[ 0 ]
  //: input g33 (B) @(80,131) /sn:0 /w:[ 0 ]
  //: input g30 (C) @(35,146) /sn:0 /w:[ 0 ]

endmodule
